library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity my_rom is
  port(
    clk : in std_logic;
    addr : in std_logic_vector(15 downto 0); -- 16 words total
    data : out std_logic_vector(5 downto 0) -- 6-bit words, RRGGBB
  );
end;

architecture sim of my_rom is
begin
  process(clk) begin
    if rising_edge(clk) then
      case addr is
        when "0000000000000000" => data <= "110000";
        when "0000000000000001" => data <= "110000";
        when "0000000000000010" => data <= "110000";
        when "0000000000000011" => data <= "110000";
        when "0000000000000100" => data <= "110000";
        when "0000000000000101" => data <= "110000";
        when "0000000000000110" => data <= "110000";
        when "0000000000000111" => data <= "110000";
        when "0000000000001000" => data <= "110000";
        when "0000000000001001" => data <= "110000";
        when "0000000000001010" => data <= "110000";
        when "0000000000001011" => data <= "110000";
        when "0000000000001100" => data <= "110000";
        when "0000000000001101" => data <= "110000";
        when "0000000000001110" => data <= "110000";
        when "0000000000001111" => data <= "110000";
        when "0000000000010000" => data <= "110000";
        when "0000000000010001" => data <= "110000";
        when "0000000000010010" => data <= "110000";
        when "0000000000010011" => data <= "110000";
        when "0000000000010100" => data <= "110000";
        when "0000000000010101" => data <= "110000";
        when "0000000000010110" => data <= "110000";
        when "0000000000010111" => data <= "110000";
        when "0000000000011000" => data <= "110000";
        when "0000000000011001" => data <= "110000";
        when "0000000000011010" => data <= "110000";
        when "0000000000011011" => data <= "110000";
        when "0000000000011100" => data <= "110000";
        when "0000000000011101" => data <= "110000";
        when "0000000000011110" => data <= "110000";
        when "0000000000011111" => data <= "110000";
        when "0000000000100000" => data <= "110000";
        when "0000000000100001" => data <= "110000";
        when "0000000000100010" => data <= "110000";
        when "0000000000100011" => data <= "110000";
        when "0000000000100100" => data <= "110000";
        when "0000000000100101" => data <= "110000";
        when "0000000000100110" => data <= "110000";
        when "0000000000100111" => data <= "110000";
        when "0000000000101000" => data <= "110000";
        when "0000000000101001" => data <= "110000";
        when "0000000000101010" => data <= "110000";
        when "0000000000101011" => data <= "110000";
        when "0000000000101100" => data <= "110000";
        when "0000000000101101" => data <= "110000";
        when "0000000000101110" => data <= "110000";
        when "0000000000101111" => data <= "110000";
        when "0000000000110000" => data <= "110000";
        when "0000000000110001" => data <= "110000";
        when "0000000000110010" => data <= "110000";
        when "0000000000110011" => data <= "110000";
        when "0000000000110100" => data <= "110000";
        when "0000000000110101" => data <= "110000";
        when "0000000000110110" => data <= "110000";
        when "0000000000110111" => data <= "110000";
        when "0000000000111000" => data <= "110000";
        when "0000000000111001" => data <= "110000";
        when "0000000000111010" => data <= "110000";
        when "0000000000111011" => data <= "110000";
        when "0000000000111100" => data <= "110000";
        when "0000000000111101" => data <= "110000";
        when "0000000000111110" => data <= "110000";
        when "0000000000111111" => data <= "110000";
        when "0000000001000000" => data <= "110000";
        when "0000000001000001" => data <= "110000";
        when "0000000001000010" => data <= "110000";
        when "0000000001000011" => data <= "110000";
        when "0000000001000100" => data <= "110000";
        when "0000000001000101" => data <= "110000";
        when "0000000001000110" => data <= "110000";
        when "0000000001000111" => data <= "110000";
        when "0000000001001000" => data <= "110000";
        when "0000000001001001" => data <= "110000";
        when "0000000001001010" => data <= "110000";
        when "0000000001001011" => data <= "110000";
        when "0000000001001100" => data <= "110000";
        when "0000000001001101" => data <= "110000";
        when "0000000001001110" => data <= "110000";
        when "0000000001001111" => data <= "110000";
        when "0000000001010000" => data <= "110000";
        when "0000000001010001" => data <= "110000";
        when "0000000001010010" => data <= "110000";
        when "0000000001010011" => data <= "110000";
        when "0000000001010100" => data <= "110000";
        when "0000000001010101" => data <= "110000";
        when "0000000001010110" => data <= "110000";
        when "0000000001010111" => data <= "110000";
        when "0000000001011000" => data <= "110000";
        when "0000000001011001" => data <= "110000";
        when "0000000001011010" => data <= "110000";
        when "0000000001011011" => data <= "110000";
        when "0000000001011100" => data <= "110000";
        when "0000000001011101" => data <= "110000";
        when "0000000001011110" => data <= "110000";
        when "0000000001011111" => data <= "110000";
        when "0000000001100000" => data <= "110000";
        when "0000000001100001" => data <= "110000";
        when "0000000001100010" => data <= "110000";
        when "0000000001100011" => data <= "110000";
        when "0000000001100100" => data <= "110000";
        when "0000000001100101" => data <= "110000";
        when "0000000001100110" => data <= "110000";
        when "0000000001100111" => data <= "110000";
        when "0000000001101000" => data <= "110000";
        when "0000000001101001" => data <= "110000";
        when "0000000001101010" => data <= "110000";
        when "0000000001101011" => data <= "110000";
        when "0000000001101100" => data <= "110000";
        when "0000000001101101" => data <= "110000";
        when "0000000001101110" => data <= "110000";
        when "0000000001101111" => data <= "110000";
        when "0000000001110000" => data <= "110000";
        when "0000000001110001" => data <= "110000";
        when "0000000001110010" => data <= "110000";
        when "0000000001110011" => data <= "110000";
        when "0000000001110100" => data <= "110000";
        when "0000000001110101" => data <= "110000";
        when "0000000001110110" => data <= "110000";
        when "0000000001110111" => data <= "110000";
        when "0000000001111000" => data <= "110000";
        when "0000000001111001" => data <= "110000";
        when "0000000001111010" => data <= "110000";
        when "0000000001111011" => data <= "110000";
        when "0000000001111100" => data <= "110000";
        when "0000000001111101" => data <= "110000";
        when "0000000001111110" => data <= "110000";
        when "0000000001111111" => data <= "110000";
        when "0000000010000000" => data <= "110000";
        when "0000000010000001" => data <= "110000";
        when "0000000010000010" => data <= "110000";
        when "0000000010000011" => data <= "110000";
        when "0000000010000100" => data <= "110000";
        when "0000000010000101" => data <= "110000";
        when "0000000010000110" => data <= "110000";
        when "0000000010000111" => data <= "110000";
        when "0000000010001000" => data <= "110000";
        when "0000000010001001" => data <= "110000";
        when "0000000010001010" => data <= "110000";
        when "0000000010001011" => data <= "110000";
        when "0000000010001100" => data <= "110000";
        when "0000000010001101" => data <= "110000";
        when "0000000010001110" => data <= "110000";
        when "0000000010001111" => data <= "110000";
        when "0000000010010000" => data <= "110000";
        when "0000000010010001" => data <= "110000";
        when "0000000010010010" => data <= "110000";
        when "0000000010010011" => data <= "110000";
        when "0000000010010100" => data <= "110000";
        when "0000000010010101" => data <= "110000";
        when "0000000010010110" => data <= "110000";
        when "0000000010010111" => data <= "110000";
        when "0000000010011000" => data <= "110000";
        when "0000000010011001" => data <= "110000";
        when "0000000010011010" => data <= "110000";
        when "0000000010011011" => data <= "110000";
        when "0000000010011100" => data <= "110000";
        when "0000000010011101" => data <= "110000";
        when "0000000010011110" => data <= "110000";
        when "0000000010011111" => data <= "110000";
        when "0000000100000000" => data <= "110000";
        when "0000000100000001" => data <= "110000";
        when "0000000100000010" => data <= "110000";
        when "0000000100000011" => data <= "110000";
        when "0000000100000100" => data <= "110000";
        when "0000000100000101" => data <= "110000";
        when "0000000100000110" => data <= "110000";
        when "0000000100000111" => data <= "110000";
        when "0000000100001000" => data <= "110000";
        when "0000000100001001" => data <= "110000";
        when "0000000100001010" => data <= "110000";
        when "0000000100001011" => data <= "110000";
        when "0000000100001100" => data <= "110000";
        when "0000000100001101" => data <= "110000";
        when "0000000100001110" => data <= "110000";
        when "0000000100001111" => data <= "110000";
        when "0000000100010000" => data <= "110000";
        when "0000000100010001" => data <= "110000";
        when "0000000100010010" => data <= "110000";
        when "0000000100010011" => data <= "110000";
        when "0000000100010100" => data <= "110000";
        when "0000000100010101" => data <= "110000";
        when "0000000100010110" => data <= "110000";
        when "0000000100010111" => data <= "110000";
        when "0000000100011000" => data <= "110000";
        when "0000000100011001" => data <= "110000";
        when "0000000100011010" => data <= "110000";
        when "0000000100011011" => data <= "110000";
        when "0000000100011100" => data <= "110000";
        when "0000000100011101" => data <= "110000";
        when "0000000100011110" => data <= "110000";
        when "0000000100011111" => data <= "110000";
        when "0000000100100000" => data <= "110000";
        when "0000000100100001" => data <= "110000";
        when "0000000100100010" => data <= "110000";
        when "0000000100100011" => data <= "110000";
        when "0000000100100100" => data <= "110000";
        when "0000000100100101" => data <= "110000";
        when "0000000100100110" => data <= "110000";
        when "0000000100100111" => data <= "110000";
        when "0000000100101000" => data <= "110000";
        when "0000000100101001" => data <= "110000";
        when "0000000100101010" => data <= "110000";
        when "0000000100101011" => data <= "110000";
        when "0000000100101100" => data <= "110000";
        when "0000000100101101" => data <= "110000";
        when "0000000100101110" => data <= "110000";
        when "0000000100101111" => data <= "110000";
        when "0000000100110000" => data <= "110000";
        when "0000000100110001" => data <= "110000";
        when "0000000100110010" => data <= "110000";
        when "0000000100110011" => data <= "110000";
        when "0000000100110100" => data <= "110000";
        when "0000000100110101" => data <= "110000";
        when "0000000100110110" => data <= "110000";
        when "0000000100110111" => data <= "110000";
        when "0000000100111000" => data <= "110000";
        when "0000000100111001" => data <= "110000";
        when "0000000100111010" => data <= "110000";
        when "0000000100111011" => data <= "110000";
        when "0000000100111100" => data <= "110000";
        when "0000000100111101" => data <= "110000";
        when "0000000100111110" => data <= "110000";
        when "0000000100111111" => data <= "110000";
        when "0000000101000000" => data <= "110000";
        when "0000000101000001" => data <= "110000";
        when "0000000101000010" => data <= "110000";
        when "0000000101000011" => data <= "110000";
        when "0000000101000100" => data <= "110000";
        when "0000000101000101" => data <= "110000";
        when "0000000101000110" => data <= "110000";
        when "0000000101000111" => data <= "110000";
        when "0000000101001000" => data <= "110000";
        when "0000000101001001" => data <= "110000";
        when "0000000101001010" => data <= "110000";
        when "0000000101001011" => data <= "110000";
        when "0000000101001100" => data <= "110000";
        when "0000000101001101" => data <= "110000";
        when "0000000101001110" => data <= "110000";
        when "0000000101001111" => data <= "110000";
        when "0000000101010000" => data <= "110000";
        when "0000000101010001" => data <= "110000";
        when "0000000101010010" => data <= "110000";
        when "0000000101010011" => data <= "110000";
        when "0000000101010100" => data <= "110000";
        when "0000000101010101" => data <= "110000";
        when "0000000101010110" => data <= "110000";
        when "0000000101010111" => data <= "110000";
        when "0000000101011000" => data <= "110000";
        when "0000000101011001" => data <= "110000";
        when "0000000101011010" => data <= "110000";
        when "0000000101011011" => data <= "110000";
        when "0000000101011100" => data <= "110000";
        when "0000000101011101" => data <= "110000";
        when "0000000101011110" => data <= "110000";
        when "0000000101011111" => data <= "110000";
        when "0000000101100000" => data <= "110000";
        when "0000000101100001" => data <= "110000";
        when "0000000101100010" => data <= "110000";
        when "0000000101100011" => data <= "110000";
        when "0000000101100100" => data <= "110000";
        when "0000000101100101" => data <= "110000";
        when "0000000101100110" => data <= "110000";
        when "0000000101100111" => data <= "110000";
        when "0000000101101000" => data <= "110000";
        when "0000000101101001" => data <= "110000";
        when "0000000101101010" => data <= "110000";
        when "0000000101101011" => data <= "110000";
        when "0000000101101100" => data <= "110000";
        when "0000000101101101" => data <= "110000";
        when "0000000101101110" => data <= "110000";
        when "0000000101101111" => data <= "110000";
        when "0000000101110000" => data <= "110000";
        when "0000000101110001" => data <= "110000";
        when "0000000101110010" => data <= "110000";
        when "0000000101110011" => data <= "110000";
        when "0000000101110100" => data <= "110000";
        when "0000000101110101" => data <= "110000";
        when "0000000101110110" => data <= "110000";
        when "0000000101110111" => data <= "110000";
        when "0000000101111000" => data <= "110000";
        when "0000000101111001" => data <= "110000";
        when "0000000101111010" => data <= "110000";
        when "0000000101111011" => data <= "110000";
        when "0000000101111100" => data <= "110000";
        when "0000000101111101" => data <= "110000";
        when "0000000101111110" => data <= "110000";
        when "0000000101111111" => data <= "110000";
        when "0000000110000000" => data <= "110000";
        when "0000000110000001" => data <= "110000";
        when "0000000110000010" => data <= "110000";
        when "0000000110000011" => data <= "110000";
        when "0000000110000100" => data <= "110000";
        when "0000000110000101" => data <= "110000";
        when "0000000110000110" => data <= "110000";
        when "0000000110000111" => data <= "110000";
        when "0000000110001000" => data <= "110000";
        when "0000000110001001" => data <= "110000";
        when "0000000110001010" => data <= "110000";
        when "0000000110001011" => data <= "110000";
        when "0000000110001100" => data <= "110000";
        when "0000000110001101" => data <= "110000";
        when "0000000110001110" => data <= "110000";
        when "0000000110001111" => data <= "110000";
        when "0000000110010000" => data <= "110000";
        when "0000000110010001" => data <= "110000";
        when "0000000110010010" => data <= "110000";
        when "0000000110010011" => data <= "110000";
        when "0000000110010100" => data <= "110000";
        when "0000000110010101" => data <= "110000";
        when "0000000110010110" => data <= "110000";
        when "0000000110010111" => data <= "110000";
        when "0000000110011000" => data <= "110000";
        when "0000000110011001" => data <= "110000";
        when "0000000110011010" => data <= "110000";
        when "0000000110011011" => data <= "110000";
        when "0000000110011100" => data <= "110000";
        when "0000000110011101" => data <= "110000";
        when "0000000110011110" => data <= "110000";
        when "0000000110011111" => data <= "110000";
        when "0000001000000000" => data <= "110000";
        when "0000001000000001" => data <= "110000";
        when "0000001001001010" => data <= "110000";
        when "0000001001001011" => data <= "110000";
        when "0000001001001100" => data <= "001001";
        when "0000001001001101" => data <= "110000";
        when "0000001001010011" => data <= "110000";
        when "0000001001010100" => data <= "110000";
        when "0000001001010101" => data <= "110000";
        when "0000001001010110" => data <= "110000";
        when "0000001010011110" => data <= "110000";
        when "0000001010011111" => data <= "110000";
        when "0000001100000000" => data <= "110000";
        when "0000001100000001" => data <= "110000";
        when "0000001100001000" => data <= "111111";
        when "0000001100001100" => data <= "111111";
        when "0000001100010000" => data <= "111111";
        when "0000001101001000" => data <= "110000";
        when "0000001101001001" => data <= "110000";
        when "0000001101001010" => data <= "001001";
        when "0000001101001011" => data <= "001001";
        when "0000001101001100" => data <= "110000";
        when "0000001101010100" => data <= "110000";
        when "0000001101010101" => data <= "001001";
        when "0000001101010110" => data <= "001001";
        when "0000001101010111" => data <= "110000";
        when "0000001101011000" => data <= "110000";
        when "0000001110001111" => data <= "111111";
        when "0000001110010011" => data <= "111111";
        when "0000001110010111" => data <= "111111";
        when "0000001110011110" => data <= "110000";
        when "0000001110011111" => data <= "110000";
        when "0000010000000000" => data <= "110000";
        when "0000010000000001" => data <= "110000";
        when "0000010000001001" => data <= "111111";
        when "0000010000001100" => data <= "111111";
        when "0000010000001111" => data <= "111111";
        when "0000010001000110" => data <= "110000";
        when "0000010001000111" => data <= "110000";
        when "0000010001001000" => data <= "001001";
        when "0000010001001001" => data <= "001001";
        when "0000010001001010" => data <= "110000";
        when "0000010001001011" => data <= "110000";
        when "0000010001010101" => data <= "110000";
        when "0000010001010110" => data <= "110000";
        when "0000010001010111" => data <= "001001";
        when "0000010001011000" => data <= "001001";
        when "0000010001011001" => data <= "110000";
        when "0000010001011010" => data <= "110000";
        when "0000010010010000" => data <= "111111";
        when "0000010010010011" => data <= "111111";
        when "0000010010010110" => data <= "111111";
        when "0000010010011110" => data <= "110000";
        when "0000010010011111" => data <= "110000";
        when "0000010100000000" => data <= "110000";
        when "0000010100000001" => data <= "110000";
        when "0000010100001010" => data <= "111111";
        when "0000010100001100" => data <= "111111";
        when "0000010100001110" => data <= "111111";
        when "0000010101000011" => data <= "110000";
        when "0000010101000100" => data <= "110000";
        when "0000010101000101" => data <= "110000";
        when "0000010101000110" => data <= "001001";
        when "0000010101000111" => data <= "001001";
        when "0000010101001000" => data <= "001001";
        when "0000010101001001" => data <= "110000";
        when "0000010101010111" => data <= "110000";
        when "0000010101011000" => data <= "001001";
        when "0000010101011001" => data <= "001001";
        when "0000010101011010" => data <= "001001";
        when "0000010101011011" => data <= "110000";
        when "0000010101011100" => data <= "110000";
        when "0000010110010001" => data <= "111111";
        when "0000010110010011" => data <= "111111";
        when "0000010110010101" => data <= "111111";
        when "0000010110011110" => data <= "110000";
        when "0000010110011111" => data <= "110000";
        when "0000011000000000" => data <= "110000";
        when "0000011000000001" => data <= "110000";
        when "0000011000001000" => data <= "111111";
        when "0000011000001011" => data <= "111111";
        when "0000011000001100" => data <= "111111";
        when "0000011000001101" => data <= "111111";
        when "0000011000010000" => data <= "111111";
        when "0000011001000001" => data <= "110000";
        when "0000011001000010" => data <= "110000";
        when "0000011001000011" => data <= "001001";
        when "0000011001000100" => data <= "001001";
        when "0000011001000101" => data <= "001001";
        when "0000011001000110" => data <= "001001";
        when "0000011001000111" => data <= "001001";
        when "0000011001001000" => data <= "110000";
        when "0000011001011000" => data <= "110000";
        when "0000011001011001" => data <= "001001";
        when "0000011001011010" => data <= "001001";
        when "0000011001011011" => data <= "001001";
        when "0000011001011100" => data <= "001001";
        when "0000011001011101" => data <= "110000";
        when "0000011001011110" => data <= "110000";
        when "0000011001011111" => data <= "110000";
        when "0000011010001111" => data <= "111111";
        when "0000011010010010" => data <= "111111";
        when "0000011010010011" => data <= "111111";
        when "0000011010010100" => data <= "111111";
        when "0000011010010111" => data <= "111111";
        when "0000011010011110" => data <= "110000";
        when "0000011010011111" => data <= "110000";
        when "0000011100000000" => data <= "110000";
        when "0000011100000001" => data <= "110000";
        when "0000011100000110" => data <= "111111";
        when "0000011100001000" => data <= "111111";
        when "0000011100001100" => data <= "111111";
        when "0000011100010000" => data <= "111111";
        when "0000011100010010" => data <= "111111";
        when "0000011100111111" => data <= "110000";
        when "0000011101000000" => data <= "110000";
        when "0000011101000001" => data <= "001001";
        when "0000011101000010" => data <= "001001";
        when "0000011101000011" => data <= "001001";
        when "0000011101000100" => data <= "001001";
        when "0000011101000101" => data <= "001001";
        when "0000011101000110" => data <= "110000";
        when "0000011101000111" => data <= "110000";
        when "0000011101011001" => data <= "110000";
        when "0000011101011010" => data <= "110000";
        when "0000011101011011" => data <= "001001";
        when "0000011101011100" => data <= "001001";
        when "0000011101011101" => data <= "001001";
        when "0000011101011110" => data <= "001001";
        when "0000011101011111" => data <= "001001";
        when "0000011101100000" => data <= "110000";
        when "0000011101100001" => data <= "110000";
        when "0000011110001101" => data <= "111111";
        when "0000011110001111" => data <= "111111";
        when "0000011110010011" => data <= "111111";
        when "0000011110010111" => data <= "111111";
        when "0000011110011001" => data <= "111111";
        when "0000011110011110" => data <= "110000";
        when "0000011110011111" => data <= "110000";
        when "0000100000000000" => data <= "110000";
        when "0000100000000001" => data <= "110000";
        when "0000100000000111" => data <= "111111";
        when "0000100000001000" => data <= "111111";
        when "0000100000001100" => data <= "111111";
        when "0000100000010000" => data <= "111111";
        when "0000100000010001" => data <= "111111";
        when "0000100000111101" => data <= "110000";
        when "0000100000111110" => data <= "110000";
        when "0000100000111111" => data <= "001001";
        when "0000100001000000" => data <= "001001";
        when "0000100001000001" => data <= "001001";
        when "0000100001000010" => data <= "001001";
        when "0000100001000011" => data <= "001001";
        when "0000100001000100" => data <= "001001";
        when "0000100001000101" => data <= "110000";
        when "0000100001011011" => data <= "110000";
        when "0000100001011100" => data <= "001001";
        when "0000100001011101" => data <= "001001";
        when "0000100001011110" => data <= "001001";
        when "0000100001011111" => data <= "001001";
        when "0000100001100000" => data <= "001001";
        when "0000100001100001" => data <= "001001";
        when "0000100001100010" => data <= "110000";
        when "0000100001100011" => data <= "110000";
        when "0000100010001110" => data <= "111111";
        when "0000100010001111" => data <= "111111";
        when "0000100010010011" => data <= "111111";
        when "0000100010010111" => data <= "111111";
        when "0000100010011000" => data <= "111111";
        when "0000100010011110" => data <= "110000";
        when "0000100010011111" => data <= "110000";
        when "0000100100000000" => data <= "110000";
        when "0000100100000001" => data <= "110000";
        when "0000100100000100" => data <= "111111";
        when "0000100100000101" => data <= "111111";
        when "0000100100000110" => data <= "111111";
        when "0000100100000111" => data <= "111111";
        when "0000100100001000" => data <= "111111";
        when "0000100100001100" => data <= "111111";
        when "0000100100010000" => data <= "111111";
        when "0000100100010001" => data <= "111111";
        when "0000100100010010" => data <= "111111";
        when "0000100100010011" => data <= "111111";
        when "0000100100010100" => data <= "111111";
        when "0000100100111010" => data <= "110000";
        when "0000100100111011" => data <= "110000";
        when "0000100100111100" => data <= "110000";
        when "0000100100111101" => data <= "001001";
        when "0000100100111110" => data <= "001001";
        when "0000100100111111" => data <= "001001";
        when "0000100101000000" => data <= "001001";
        when "0000100101000001" => data <= "001001";
        when "0000100101000010" => data <= "001001";
        when "0000100101000011" => data <= "001001";
        when "0000100101000100" => data <= "110000";
        when "0000100101001001" => data <= "110000";
        when "0000100101001010" => data <= "110000";
        when "0000100101001011" => data <= "110000";
        when "0000100101001100" => data <= "110000";
        when "0000100101001101" => data <= "110000";
        when "0000100101001110" => data <= "110000";
        when "0000100101001111" => data <= "110000";
        when "0000100101010000" => data <= "110000";
        when "0000100101010001" => data <= "110000";
        when "0000100101010010" => data <= "110000";
        when "0000100101010011" => data <= "110000";
        when "0000100101010100" => data <= "110000";
        when "0000100101010101" => data <= "110000";
        when "0000100101010110" => data <= "110000";
        when "0000100101010111" => data <= "110000";
        when "0000100101011100" => data <= "110000";
        when "0000100101011101" => data <= "001001";
        when "0000100101011110" => data <= "001001";
        when "0000100101011111" => data <= "001001";
        when "0000100101100000" => data <= "001001";
        when "0000100101100001" => data <= "001001";
        when "0000100101100010" => data <= "001001";
        when "0000100101100011" => data <= "001001";
        when "0000100101100100" => data <= "110000";
        when "0000100101100101" => data <= "110000";
        when "0000100110001011" => data <= "111111";
        when "0000100110001100" => data <= "111111";
        when "0000100110001101" => data <= "111111";
        when "0000100110001110" => data <= "111111";
        when "0000100110001111" => data <= "111111";
        when "0000100110010011" => data <= "111111";
        when "0000100110010111" => data <= "111111";
        when "0000100110011000" => data <= "111111";
        when "0000100110011001" => data <= "111111";
        when "0000100110011010" => data <= "111111";
        when "0000100110011011" => data <= "111111";
        when "0000100110011110" => data <= "110000";
        when "0000100110011111" => data <= "110000";
        when "0000101000000000" => data <= "110000";
        when "0000101000000001" => data <= "110000";
        when "0000101000001001" => data <= "111111";
        when "0000101000001100" => data <= "111111";
        when "0000101000001111" => data <= "111111";
        when "0000101000111000" => data <= "110000";
        when "0000101000111001" => data <= "110000";
        when "0000101000111010" => data <= "001001";
        when "0000101000111011" => data <= "001001";
        when "0000101000111100" => data <= "001001";
        when "0000101000111101" => data <= "001001";
        when "0000101000111110" => data <= "001001";
        when "0000101000111111" => data <= "001001";
        when "0000101001000000" => data <= "001001";
        when "0000101001000001" => data <= "001001";
        when "0000101001000010" => data <= "110000";
        when "0000101001000011" => data <= "110000";
        when "0000101001001001" => data <= "110000";
        when "0000101001010111" => data <= "110000";
        when "0000101001011101" => data <= "110000";
        when "0000101001011110" => data <= "110000";
        when "0000101001011111" => data <= "001001";
        when "0000101001100000" => data <= "001001";
        when "0000101001100001" => data <= "001001";
        when "0000101001100010" => data <= "001001";
        when "0000101001100011" => data <= "001001";
        when "0000101001100100" => data <= "001001";
        when "0000101001100101" => data <= "001001";
        when "0000101001100110" => data <= "110000";
        when "0000101001100111" => data <= "110000";
        when "0000101010010000" => data <= "111111";
        when "0000101010010011" => data <= "111111";
        when "0000101010010110" => data <= "111111";
        when "0000101010011110" => data <= "110000";
        when "0000101010011111" => data <= "110000";
        when "0000101100000000" => data <= "110000";
        when "0000101100000001" => data <= "110000";
        when "0000101100000101" => data <= "111111";
        when "0000101100001010" => data <= "111111";
        when "0000101100001100" => data <= "111111";
        when "0000101100001110" => data <= "111111";
        when "0000101100010011" => data <= "111111";
        when "0000101100110110" => data <= "110000";
        when "0000101100110111" => data <= "110000";
        when "0000101100111000" => data <= "001001";
        when "0000101100111001" => data <= "001001";
        when "0000101100111010" => data <= "001001";
        when "0000101100111011" => data <= "001001";
        when "0000101100111100" => data <= "001001";
        when "0000101100111101" => data <= "001001";
        when "0000101100111110" => data <= "001001";
        when "0000101100111111" => data <= "001001";
        when "0000101101000000" => data <= "001001";
        when "0000101101000001" => data <= "110000";
        when "0000101101001001" => data <= "110000";
        when "0000101101010111" => data <= "110000";
        when "0000101101011111" => data <= "110000";
        when "0000101101100000" => data <= "001001";
        when "0000101101100001" => data <= "001001";
        when "0000101101100010" => data <= "001001";
        when "0000101101100011" => data <= "001001";
        when "0000101101100100" => data <= "001001";
        when "0000101101100101" => data <= "001001";
        when "0000101101100110" => data <= "001001";
        when "0000101101100111" => data <= "001001";
        when "0000101101101000" => data <= "110000";
        when "0000101101101001" => data <= "110000";
        when "0000101101101010" => data <= "110000";
        when "0000101110001100" => data <= "111111";
        when "0000101110010001" => data <= "111111";
        when "0000101110010011" => data <= "111111";
        when "0000101110010101" => data <= "111111";
        when "0000101110011010" => data <= "111111";
        when "0000101110011110" => data <= "110000";
        when "0000101110011111" => data <= "110000";
        when "0000110000000000" => data <= "110000";
        when "0000110000000001" => data <= "110000";
        when "0000110000000110" => data <= "111111";
        when "0000110000001011" => data <= "111111";
        when "0000110000001100" => data <= "111111";
        when "0000110000001101" => data <= "111111";
        when "0000110000010010" => data <= "111111";
        when "0000110000110100" => data <= "110000";
        when "0000110000110101" => data <= "110000";
        when "0000110000110110" => data <= "001001";
        when "0000110000110111" => data <= "001001";
        when "0000110000111000" => data <= "001001";
        when "0000110000111001" => data <= "001001";
        when "0000110000111010" => data <= "001001";
        when "0000110000111011" => data <= "001001";
        when "0000110000111100" => data <= "001001";
        when "0000110000111101" => data <= "001001";
        when "0000110000111110" => data <= "001001";
        when "0000110000111111" => data <= "110000";
        when "0000110001000000" => data <= "110000";
        when "0000110001001001" => data <= "110000";
        when "0000110001010111" => data <= "110000";
        when "0000110001100000" => data <= "110000";
        when "0000110001100001" => data <= "001001";
        when "0000110001100010" => data <= "001001";
        when "0000110001100011" => data <= "001001";
        when "0000110001100100" => data <= "001001";
        when "0000110001100101" => data <= "001001";
        when "0000110001100110" => data <= "001001";
        when "0000110001100111" => data <= "001001";
        when "0000110001101000" => data <= "001001";
        when "0000110001101001" => data <= "001001";
        when "0000110001101010" => data <= "001001";
        when "0000110001101011" => data <= "110000";
        when "0000110001101100" => data <= "110000";
        when "0000110010001101" => data <= "111111";
        when "0000110010010010" => data <= "111111";
        when "0000110010010011" => data <= "111111";
        when "0000110010010100" => data <= "111111";
        when "0000110010011001" => data <= "111111";
        when "0000110010011110" => data <= "110000";
        when "0000110010011111" => data <= "110000";
        when "0000110100000000" => data <= "110000";
        when "0000110100000001" => data <= "110000";
        when "0000110100000011" => data <= "111111";
        when "0000110100000100" => data <= "111111";
        when "0000110100000101" => data <= "111111";
        when "0000110100000110" => data <= "111111";
        when "0000110100000111" => data <= "111111";
        when "0000110100001000" => data <= "111111";
        when "0000110100001001" => data <= "111111";
        when "0000110100001010" => data <= "111111";
        when "0000110100001011" => data <= "111111";
        when "0000110100001100" => data <= "111111";
        when "0000110100001101" => data <= "111111";
        when "0000110100001110" => data <= "111111";
        when "0000110100001111" => data <= "111111";
        when "0000110100010000" => data <= "111111";
        when "0000110100010001" => data <= "111111";
        when "0000110100010010" => data <= "111111";
        when "0000110100010011" => data <= "111111";
        when "0000110100010100" => data <= "111111";
        when "0000110100010101" => data <= "111111";
        when "0000110100110001" => data <= "110000";
        when "0000110100110010" => data <= "110000";
        when "0000110100110011" => data <= "110000";
        when "0000110100110100" => data <= "001001";
        when "0000110100110101" => data <= "001001";
        when "0000110100110110" => data <= "001001";
        when "0000110100110111" => data <= "001001";
        when "0000110100111000" => data <= "001001";
        when "0000110100111001" => data <= "001001";
        when "0000110100111010" => data <= "001001";
        when "0000110100111011" => data <= "001001";
        when "0000110100111100" => data <= "001001";
        when "0000110100111101" => data <= "001001";
        when "0000110100111110" => data <= "110000";
        when "0000110101001001" => data <= "110000";
        when "0000110101010111" => data <= "110000";
        when "0000110101100001" => data <= "110000";
        when "0000110101100010" => data <= "110000";
        when "0000110101100011" => data <= "001001";
        when "0000110101100100" => data <= "001001";
        when "0000110101100101" => data <= "001001";
        when "0000110101100110" => data <= "001001";
        when "0000110101100111" => data <= "001001";
        when "0000110101101000" => data <= "001001";
        when "0000110101101001" => data <= "001001";
        when "0000110101101010" => data <= "001001";
        when "0000110101101011" => data <= "001001";
        when "0000110101101100" => data <= "001001";
        when "0000110101101101" => data <= "110000";
        when "0000110101101110" => data <= "110000";
        when "0000110110001010" => data <= "111111";
        when "0000110110001011" => data <= "111111";
        when "0000110110001100" => data <= "111111";
        when "0000110110001101" => data <= "111111";
        when "0000110110001110" => data <= "111111";
        when "0000110110001111" => data <= "111111";
        when "0000110110010000" => data <= "111111";
        when "0000110110010001" => data <= "111111";
        when "0000110110010010" => data <= "111111";
        when "0000110110010011" => data <= "111111";
        when "0000110110010100" => data <= "111111";
        when "0000110110010101" => data <= "111111";
        when "0000110110010110" => data <= "111111";
        when "0000110110010111" => data <= "111111";
        when "0000110110011000" => data <= "111111";
        when "0000110110011001" => data <= "111111";
        when "0000110110011010" => data <= "111111";
        when "0000110110011011" => data <= "111111";
        when "0000110110011100" => data <= "111111";
        when "0000110110011110" => data <= "110000";
        when "0000110110011111" => data <= "110000";
        when "0000111000000000" => data <= "110000";
        when "0000111000000001" => data <= "110000";
        when "0000111000000110" => data <= "111111";
        when "0000111000001011" => data <= "111111";
        when "0000111000001100" => data <= "111111";
        when "0000111000001101" => data <= "111111";
        when "0000111000010010" => data <= "111111";
        when "0000111000101111" => data <= "110000";
        when "0000111000110000" => data <= "110000";
        when "0000111000110001" => data <= "001001";
        when "0000111000110010" => data <= "001001";
        when "0000111000110011" => data <= "001001";
        when "0000111000110100" => data <= "001001";
        when "0000111000110101" => data <= "001001";
        when "0000111000110110" => data <= "001001";
        when "0000111000110111" => data <= "001001";
        when "0000111000111000" => data <= "001001";
        when "0000111000111001" => data <= "001001";
        when "0000111000111010" => data <= "001001";
        when "0000111000111011" => data <= "001001";
        when "0000111000111100" => data <= "001001";
        when "0000111000111101" => data <= "110000";
        when "0000111001001001" => data <= "110000";
        when "0000111001010111" => data <= "110000";
        when "0000111001100011" => data <= "110000";
        when "0000111001100100" => data <= "001001";
        when "0000111001100101" => data <= "001001";
        when "0000111001100110" => data <= "001001";
        when "0000111001100111" => data <= "001001";
        when "0000111001101000" => data <= "001001";
        when "0000111001101001" => data <= "001001";
        when "0000111001101010" => data <= "001001";
        when "0000111001101011" => data <= "001001";
        when "0000111001101100" => data <= "001001";
        when "0000111001101101" => data <= "001001";
        when "0000111001101110" => data <= "001001";
        when "0000111001101111" => data <= "110000";
        when "0000111001110000" => data <= "110000";
        when "0000111010001101" => data <= "111111";
        when "0000111010010010" => data <= "111111";
        when "0000111010010011" => data <= "111111";
        when "0000111010010100" => data <= "111111";
        when "0000111010011001" => data <= "111111";
        when "0000111010011110" => data <= "110000";
        when "0000111010011111" => data <= "110000";
        when "0000111100000000" => data <= "110000";
        when "0000111100000001" => data <= "110000";
        when "0000111100000101" => data <= "111111";
        when "0000111100001010" => data <= "111111";
        when "0000111100001100" => data <= "111111";
        when "0000111100001110" => data <= "111111";
        when "0000111100010011" => data <= "111111";
        when "0000111100101101" => data <= "110000";
        when "0000111100101110" => data <= "110000";
        when "0000111100101111" => data <= "001001";
        when "0000111100110000" => data <= "001001";
        when "0000111100110001" => data <= "001001";
        when "0000111100110010" => data <= "001001";
        when "0000111100110011" => data <= "001001";
        when "0000111100110100" => data <= "001001";
        when "0000111100110101" => data <= "001001";
        when "0000111100110110" => data <= "001001";
        when "0000111100110111" => data <= "001001";
        when "0000111100111000" => data <= "001001";
        when "0000111100111001" => data <= "001001";
        when "0000111100111010" => data <= "001001";
        when "0000111100111011" => data <= "110000";
        when "0000111100111100" => data <= "110000";
        when "0000111101001001" => data <= "110000";
        when "0000111101010111" => data <= "110000";
        when "0000111101100100" => data <= "110000";
        when "0000111101100101" => data <= "001001";
        when "0000111101100110" => data <= "001001";
        when "0000111101100111" => data <= "001001";
        when "0000111101101000" => data <= "001001";
        when "0000111101101001" => data <= "001001";
        when "0000111101101010" => data <= "001001";
        when "0000111101101011" => data <= "001001";
        when "0000111101101100" => data <= "001001";
        when "0000111101101101" => data <= "001001";
        when "0000111101101110" => data <= "001001";
        when "0000111101101111" => data <= "001001";
        when "0000111101110000" => data <= "001001";
        when "0000111101110001" => data <= "110000";
        when "0000111101110010" => data <= "110000";
        when "0000111101110011" => data <= "110000";
        when "0000111110001100" => data <= "111111";
        when "0000111110010001" => data <= "111111";
        when "0000111110010011" => data <= "111111";
        when "0000111110010101" => data <= "111111";
        when "0000111110011010" => data <= "111111";
        when "0000111110011110" => data <= "110000";
        when "0000111110011111" => data <= "110000";
        when "0001000000000000" => data <= "110000";
        when "0001000000000001" => data <= "110000";
        when "0001000000001001" => data <= "111111";
        when "0001000000001100" => data <= "111111";
        when "0001000000001111" => data <= "111111";
        when "0001000000101011" => data <= "110000";
        when "0001000000101100" => data <= "110000";
        when "0001000000101101" => data <= "001001";
        when "0001000000101110" => data <= "001001";
        when "0001000000101111" => data <= "001001";
        when "0001000000110000" => data <= "001001";
        when "0001000000110001" => data <= "001001";
        when "0001000000110010" => data <= "001001";
        when "0001000000110011" => data <= "001001";
        when "0001000000110100" => data <= "001001";
        when "0001000000110101" => data <= "001001";
        when "0001000000110110" => data <= "001001";
        when "0001000000110111" => data <= "001001";
        when "0001000000111000" => data <= "001001";
        when "0001000000111001" => data <= "001001";
        when "0001000000111010" => data <= "110000";
        when "0001000001001001" => data <= "110000";
        when "0001000001010111" => data <= "110000";
        when "0001000001100101" => data <= "110000";
        when "0001000001100110" => data <= "110000";
        when "0001000001100111" => data <= "001001";
        when "0001000001101000" => data <= "001001";
        when "0001000001101001" => data <= "001001";
        when "0001000001101010" => data <= "001001";
        when "0001000001101011" => data <= "001001";
        when "0001000001101100" => data <= "001001";
        when "0001000001101101" => data <= "001001";
        when "0001000001101110" => data <= "001001";
        when "0001000001101111" => data <= "001001";
        when "0001000001110000" => data <= "001001";
        when "0001000001110001" => data <= "001001";
        when "0001000001110010" => data <= "001001";
        when "0001000001110011" => data <= "001001";
        when "0001000001110100" => data <= "110000";
        when "0001000001110101" => data <= "110000";
        when "0001000010010000" => data <= "111111";
        when "0001000010010011" => data <= "111111";
        when "0001000010010110" => data <= "111111";
        when "0001000010011110" => data <= "110000";
        when "0001000010011111" => data <= "110000";
        when "0001000100000000" => data <= "110000";
        when "0001000100000001" => data <= "110000";
        when "0001000100000100" => data <= "111111";
        when "0001000100000101" => data <= "111111";
        when "0001000100000110" => data <= "111111";
        when "0001000100000111" => data <= "111111";
        when "0001000100001000" => data <= "111111";
        when "0001000100001100" => data <= "111111";
        when "0001000100010000" => data <= "111111";
        when "0001000100010001" => data <= "111111";
        when "0001000100010010" => data <= "111111";
        when "0001000100010011" => data <= "111111";
        when "0001000100010100" => data <= "111111";
        when "0001000100101000" => data <= "110000";
        when "0001000100101001" => data <= "110000";
        when "0001000100101010" => data <= "110000";
        when "0001000100101011" => data <= "001001";
        when "0001000100101100" => data <= "001001";
        when "0001000100101101" => data <= "001001";
        when "0001000100101110" => data <= "001001";
        when "0001000100101111" => data <= "001001";
        when "0001000100110000" => data <= "001001";
        when "0001000100110001" => data <= "001001";
        when "0001000100110010" => data <= "001001";
        when "0001000100110011" => data <= "001001";
        when "0001000100110100" => data <= "001001";
        when "0001000100110101" => data <= "001001";
        when "0001000100110110" => data <= "001001";
        when "0001000100110111" => data <= "001001";
        when "0001000100111000" => data <= "001001";
        when "0001000100111001" => data <= "110000";
        when "0001000101001001" => data <= "110000";
        when "0001000101010111" => data <= "110000";
        when "0001000101100111" => data <= "110000";
        when "0001000101101000" => data <= "001001";
        when "0001000101101001" => data <= "001001";
        when "0001000101101010" => data <= "001001";
        when "0001000101101011" => data <= "001001";
        when "0001000101101100" => data <= "001001";
        when "0001000101101101" => data <= "001001";
        when "0001000101101110" => data <= "001001";
        when "0001000101101111" => data <= "001001";
        when "0001000101110000" => data <= "001001";
        when "0001000101110001" => data <= "001001";
        when "0001000101110010" => data <= "001001";
        when "0001000101110011" => data <= "001001";
        when "0001000101110100" => data <= "001001";
        when "0001000101110101" => data <= "001001";
        when "0001000101110110" => data <= "110000";
        when "0001000101110111" => data <= "110000";
        when "0001000110001011" => data <= "111111";
        when "0001000110001100" => data <= "111111";
        when "0001000110001101" => data <= "111111";
        when "0001000110001110" => data <= "111111";
        when "0001000110001111" => data <= "111111";
        when "0001000110010011" => data <= "111111";
        when "0001000110010111" => data <= "111111";
        when "0001000110011000" => data <= "111111";
        when "0001000110011001" => data <= "111111";
        when "0001000110011010" => data <= "111111";
        when "0001000110011011" => data <= "111111";
        when "0001000110011110" => data <= "110000";
        when "0001000110011111" => data <= "110000";
        when "0001001000000000" => data <= "110000";
        when "0001001000000001" => data <= "110000";
        when "0001001000000111" => data <= "111111";
        when "0001001000001000" => data <= "111111";
        when "0001001000001100" => data <= "111111";
        when "0001001000010000" => data <= "111111";
        when "0001001000010001" => data <= "111111";
        when "0001001000100110" => data <= "110000";
        when "0001001000100111" => data <= "110000";
        when "0001001000101000" => data <= "001001";
        when "0001001000101001" => data <= "001001";
        when "0001001000101010" => data <= "001001";
        when "0001001000101011" => data <= "001001";
        when "0001001000101100" => data <= "001001";
        when "0001001000101101" => data <= "001001";
        when "0001001000101110" => data <= "001001";
        when "0001001000101111" => data <= "001001";
        when "0001001000110000" => data <= "001001";
        when "0001001000110001" => data <= "001001";
        when "0001001000110010" => data <= "001001";
        when "0001001000110011" => data <= "001001";
        when "0001001000110100" => data <= "001001";
        when "0001001000110101" => data <= "001001";
        when "0001001000110110" => data <= "001001";
        when "0001001000110111" => data <= "110000";
        when "0001001000111000" => data <= "110000";
        when "0001001001000110" => data <= "110000";
        when "0001001001000111" => data <= "110000";
        when "0001001001001000" => data <= "110000";
        when "0001001001001001" => data <= "110000";
        when "0001001001010011" => data <= "110000";
        when "0001001001010100" => data <= "110000";
        when "0001001001010101" => data <= "110000";
        when "0001001001010110" => data <= "110000";
        when "0001001001010111" => data <= "110000";
        when "0001001001101000" => data <= "110000";
        when "0001001001101001" => data <= "001001";
        when "0001001001101010" => data <= "001001";
        when "0001001001101011" => data <= "001001";
        when "0001001001101100" => data <= "001001";
        when "0001001001101101" => data <= "001001";
        when "0001001001101110" => data <= "001001";
        when "0001001001101111" => data <= "001001";
        when "0001001001110000" => data <= "001001";
        when "0001001001110001" => data <= "001001";
        when "0001001001110010" => data <= "001001";
        when "0001001001110011" => data <= "001001";
        when "0001001001110100" => data <= "001001";
        when "0001001001110101" => data <= "001001";
        when "0001001001110110" => data <= "001001";
        when "0001001001110111" => data <= "001001";
        when "0001001001111000" => data <= "110000";
        when "0001001001111001" => data <= "110000";
        when "0001001010001110" => data <= "111111";
        when "0001001010001111" => data <= "111111";
        when "0001001010010011" => data <= "111111";
        when "0001001010010111" => data <= "111111";
        when "0001001010011000" => data <= "111111";
        when "0001001010011110" => data <= "110000";
        when "0001001010011111" => data <= "110000";
        when "0001001100000000" => data <= "110000";
        when "0001001100000001" => data <= "110000";
        when "0001001100000110" => data <= "111111";
        when "0001001100001000" => data <= "111111";
        when "0001001100001100" => data <= "111111";
        when "0001001100010000" => data <= "111111";
        when "0001001100010010" => data <= "111111";
        when "0001001100100100" => data <= "110000";
        when "0001001100100101" => data <= "110000";
        when "0001001100100110" => data <= "001001";
        when "0001001100100111" => data <= "001001";
        when "0001001100101000" => data <= "001001";
        when "0001001100101001" => data <= "001001";
        when "0001001100101010" => data <= "001001";
        when "0001001100101011" => data <= "001001";
        when "0001001100101100" => data <= "001001";
        when "0001001100101101" => data <= "001001";
        when "0001001100101110" => data <= "001001";
        when "0001001100101111" => data <= "001001";
        when "0001001100110000" => data <= "001001";
        when "0001001100110001" => data <= "001001";
        when "0001001100110010" => data <= "001001";
        when "0001001100110011" => data <= "001001";
        when "0001001100110100" => data <= "001001";
        when "0001001100110101" => data <= "001001";
        when "0001001100110110" => data <= "110000";
        when "0001001101000110" => data <= "110000";
        when "0001001101000111" => data <= "110000";
        when "0001001101001000" => data <= "110000";
        when "0001001101001001" => data <= "110000";
        when "0001001101010011" => data <= "110000";
        when "0001001101010100" => data <= "110000";
        when "0001001101010101" => data <= "110000";
        when "0001001101010110" => data <= "110000";
        when "0001001101010111" => data <= "110000";
        when "0001001101101001" => data <= "110000";
        when "0001001101101010" => data <= "110000";
        when "0001001101101011" => data <= "001001";
        when "0001001101101100" => data <= "001001";
        when "0001001101101101" => data <= "001001";
        when "0001001101101110" => data <= "001001";
        when "0001001101101111" => data <= "001001";
        when "0001001101110000" => data <= "001001";
        when "0001001101110001" => data <= "001001";
        when "0001001101110010" => data <= "001001";
        when "0001001101110011" => data <= "001001";
        when "0001001101110100" => data <= "001001";
        when "0001001101110101" => data <= "001001";
        when "0001001101110110" => data <= "001001";
        when "0001001101110111" => data <= "001001";
        when "0001001101111000" => data <= "001001";
        when "0001001101111001" => data <= "001001";
        when "0001001101111010" => data <= "110000";
        when "0001001101111011" => data <= "110000";
        when "0001001101111100" => data <= "110000";
        when "0001001110001101" => data <= "111111";
        when "0001001110001111" => data <= "111111";
        when "0001001110010011" => data <= "111111";
        when "0001001110010111" => data <= "111111";
        when "0001001110011001" => data <= "111111";
        when "0001001110011110" => data <= "110000";
        when "0001001110011111" => data <= "110000";
        when "0001010000000000" => data <= "110000";
        when "0001010000000001" => data <= "110000";
        when "0001010000001000" => data <= "111111";
        when "0001010000001011" => data <= "111111";
        when "0001010000001100" => data <= "111111";
        when "0001010000001101" => data <= "111111";
        when "0001010000010000" => data <= "111111";
        when "0001010000100010" => data <= "110000";
        when "0001010000100011" => data <= "110000";
        when "0001010000100100" => data <= "001001";
        when "0001010000100101" => data <= "001001";
        when "0001010000100110" => data <= "001001";
        when "0001010000100111" => data <= "001001";
        when "0001010000101000" => data <= "001001";
        when "0001010000101001" => data <= "001001";
        when "0001010000101010" => data <= "001001";
        when "0001010000101011" => data <= "001001";
        when "0001010000101100" => data <= "001001";
        when "0001010000101101" => data <= "001001";
        when "0001010000101110" => data <= "001001";
        when "0001010000101111" => data <= "001001";
        when "0001010000110000" => data <= "001001";
        when "0001010000110001" => data <= "001001";
        when "0001010000110010" => data <= "001001";
        when "0001010000110011" => data <= "001001";
        when "0001010000110100" => data <= "001001";
        when "0001010000110101" => data <= "110000";
        when "0001010001000101" => data <= "110000";
        when "0001010001000110" => data <= "110000";
        when "0001010001000111" => data <= "110000";
        when "0001010001001000" => data <= "110000";
        when "0001010001001001" => data <= "110000";
        when "0001010001010010" => data <= "110000";
        when "0001010001010011" => data <= "110000";
        when "0001010001010100" => data <= "110000";
        when "0001010001010101" => data <= "110000";
        when "0001010001010110" => data <= "110000";
        when "0001010001010111" => data <= "110000";
        when "0001010001101011" => data <= "110000";
        when "0001010001101100" => data <= "001001";
        when "0001010001101101" => data <= "001001";
        when "0001010001101110" => data <= "001001";
        when "0001010001101111" => data <= "001001";
        when "0001010001110000" => data <= "001001";
        when "0001010001110001" => data <= "001001";
        when "0001010001110010" => data <= "001001";
        when "0001010001110011" => data <= "001001";
        when "0001010001110100" => data <= "001001";
        when "0001010001110101" => data <= "001001";
        when "0001010001110110" => data <= "001001";
        when "0001010001110111" => data <= "001001";
        when "0001010001111000" => data <= "001001";
        when "0001010001111001" => data <= "001001";
        when "0001010001111010" => data <= "001001";
        when "0001010001111011" => data <= "001001";
        when "0001010001111100" => data <= "001001";
        when "0001010001111101" => data <= "110000";
        when "0001010001111110" => data <= "110000";
        when "0001010010001111" => data <= "111111";
        when "0001010010010010" => data <= "111111";
        when "0001010010010011" => data <= "111111";
        when "0001010010010100" => data <= "111111";
        when "0001010010010111" => data <= "111111";
        when "0001010010011110" => data <= "110000";
        when "0001010010011111" => data <= "110000";
        when "0001010100000000" => data <= "110000";
        when "0001010100000001" => data <= "110000";
        when "0001010100001010" => data <= "111111";
        when "0001010100001100" => data <= "111111";
        when "0001010100001110" => data <= "111111";
        when "0001010100011111" => data <= "110000";
        when "0001010100100000" => data <= "110000";
        when "0001010100100001" => data <= "110000";
        when "0001010100100010" => data <= "001001";
        when "0001010100100011" => data <= "001001";
        when "0001010100100100" => data <= "001001";
        when "0001010100100101" => data <= "001001";
        when "0001010100100110" => data <= "001001";
        when "0001010100100111" => data <= "001001";
        when "0001010100101000" => data <= "001001";
        when "0001010100101001" => data <= "001001";
        when "0001010100101010" => data <= "001001";
        when "0001010100101011" => data <= "001001";
        when "0001010100101100" => data <= "001001";
        when "0001010100101101" => data <= "001001";
        when "0001010100101110" => data <= "001001";
        when "0001010100101111" => data <= "001001";
        when "0001010100110000" => data <= "001001";
        when "0001010100110001" => data <= "001001";
        when "0001010100110010" => data <= "001001";
        when "0001010100110011" => data <= "110000";
        when "0001010100110100" => data <= "110000";
        when "0001010101000101" => data <= "110000";
        when "0001010101000110" => data <= "110000";
        when "0001010101000111" => data <= "110000";
        when "0001010101001000" => data <= "110000";
        when "0001010101001001" => data <= "110000";
        when "0001010101010010" => data <= "110000";
        when "0001010101010011" => data <= "110000";
        when "0001010101010100" => data <= "110000";
        when "0001010101010101" => data <= "110000";
        when "0001010101010110" => data <= "110000";
        when "0001010101010111" => data <= "110000";
        when "0001010101101100" => data <= "110000";
        when "0001010101101101" => data <= "001001";
        when "0001010101101110" => data <= "001001";
        when "0001010101101111" => data <= "001001";
        when "0001010101110000" => data <= "001001";
        when "0001010101110001" => data <= "001001";
        when "0001010101110010" => data <= "001001";
        when "0001010101110011" => data <= "001001";
        when "0001010101110100" => data <= "001001";
        when "0001010101110101" => data <= "001001";
        when "0001010101110110" => data <= "001001";
        when "0001010101110111" => data <= "001001";
        when "0001010101111000" => data <= "001001";
        when "0001010101111001" => data <= "001001";
        when "0001010101111010" => data <= "001001";
        when "0001010101111011" => data <= "001001";
        when "0001010101111100" => data <= "001001";
        when "0001010101111101" => data <= "001001";
        when "0001010101111110" => data <= "001001";
        when "0001010101111111" => data <= "110000";
        when "0001010110000000" => data <= "110000";
        when "0001010110010001" => data <= "111111";
        when "0001010110010011" => data <= "111111";
        when "0001010110010101" => data <= "111111";
        when "0001010110011110" => data <= "110000";
        when "0001010110011111" => data <= "110000";
        when "0001011000000000" => data <= "110000";
        when "0001011000000001" => data <= "110000";
        when "0001011000001001" => data <= "111111";
        when "0001011000001100" => data <= "111111";
        when "0001011000001111" => data <= "111111";
        when "0001011000011101" => data <= "110000";
        when "0001011000011110" => data <= "110000";
        when "0001011000011111" => data <= "001001";
        when "0001011000100000" => data <= "001001";
        when "0001011000100001" => data <= "001001";
        when "0001011000100010" => data <= "001001";
        when "0001011000100011" => data <= "001001";
        when "0001011000100100" => data <= "001001";
        when "0001011000100101" => data <= "001001";
        when "0001011000100110" => data <= "001001";
        when "0001011000100111" => data <= "001001";
        when "0001011000101000" => data <= "001001";
        when "0001011000101001" => data <= "001001";
        when "0001011000101010" => data <= "001001";
        when "0001011000101011" => data <= "001001";
        when "0001011000101100" => data <= "001001";
        when "0001011000101101" => data <= "001001";
        when "0001011000101110" => data <= "001001";
        when "0001011000101111" => data <= "001001";
        when "0001011000110000" => data <= "001001";
        when "0001011000110001" => data <= "001001";
        when "0001011000110010" => data <= "110000";
        when "0001011001000101" => data <= "110000";
        when "0001011001000110" => data <= "110000";
        when "0001011001000111" => data <= "110000";
        when "0001011001001000" => data <= "110000";
        when "0001011001001001" => data <= "110000";
        when "0001011001010010" => data <= "110000";
        when "0001011001010011" => data <= "110000";
        when "0001011001010100" => data <= "110000";
        when "0001011001010101" => data <= "110000";
        when "0001011001010110" => data <= "110000";
        when "0001011001010111" => data <= "110000";
        when "0001011001101101" => data <= "110000";
        when "0001011001101110" => data <= "110000";
        when "0001011001101111" => data <= "001001";
        when "0001011001110000" => data <= "001001";
        when "0001011001110001" => data <= "001001";
        when "0001011001110010" => data <= "001001";
        when "0001011001110011" => data <= "001001";
        when "0001011001110100" => data <= "001001";
        when "0001011001110101" => data <= "001001";
        when "0001011001110110" => data <= "001001";
        when "0001011001110111" => data <= "001001";
        when "0001011001111000" => data <= "001001";
        when "0001011001111001" => data <= "001001";
        when "0001011001111010" => data <= "001001";
        when "0001011001111011" => data <= "001001";
        when "0001011001111100" => data <= "001001";
        when "0001011001111101" => data <= "001001";
        when "0001011001111110" => data <= "001001";
        when "0001011001111111" => data <= "001001";
        when "0001011010000000" => data <= "001001";
        when "0001011010000001" => data <= "110000";
        when "0001011010000010" => data <= "110000";
        when "0001011010010000" => data <= "111111";
        when "0001011010010011" => data <= "111111";
        when "0001011010010110" => data <= "111111";
        when "0001011010011110" => data <= "110000";
        when "0001011010011111" => data <= "110000";
        when "0001011100000000" => data <= "110000";
        when "0001011100000001" => data <= "110000";
        when "0001011100001000" => data <= "111111";
        when "0001011100001100" => data <= "111111";
        when "0001011100010000" => data <= "111111";
        when "0001011100011011" => data <= "110000";
        when "0001011100011100" => data <= "110000";
        when "0001011100011101" => data <= "001001";
        when "0001011100011110" => data <= "001001";
        when "0001011100011111" => data <= "001001";
        when "0001011100100000" => data <= "001001";
        when "0001011100100001" => data <= "001001";
        when "0001011100100010" => data <= "001001";
        when "0001011100100011" => data <= "001001";
        when "0001011100100100" => data <= "001001";
        when "0001011100100101" => data <= "001001";
        when "0001011100100110" => data <= "001001";
        when "0001011100100111" => data <= "001001";
        when "0001011100101000" => data <= "001001";
        when "0001011100101001" => data <= "001001";
        when "0001011100101010" => data <= "001001";
        when "0001011100101011" => data <= "001001";
        when "0001011100101100" => data <= "001001";
        when "0001011100101101" => data <= "001001";
        when "0001011100101110" => data <= "001001";
        when "0001011100101111" => data <= "001001";
        when "0001011100110000" => data <= "001001";
        when "0001011100110001" => data <= "110000";
        when "0001011101000101" => data <= "110000";
        when "0001011101000110" => data <= "110000";
        when "0001011101000111" => data <= "110000";
        when "0001011101001000" => data <= "110000";
        when "0001011101001001" => data <= "110000";
        when "0001011101010010" => data <= "110000";
        when "0001011101010011" => data <= "110000";
        when "0001011101010100" => data <= "110000";
        when "0001011101010101" => data <= "110000";
        when "0001011101010110" => data <= "110000";
        when "0001011101010111" => data <= "110000";
        when "0001011101101111" => data <= "110000";
        when "0001011101110000" => data <= "001001";
        when "0001011101110001" => data <= "001001";
        when "0001011101110010" => data <= "001001";
        when "0001011101110011" => data <= "001001";
        when "0001011101110100" => data <= "001001";
        when "0001011101110101" => data <= "001001";
        when "0001011101110110" => data <= "001001";
        when "0001011101110111" => data <= "001001";
        when "0001011101111000" => data <= "001001";
        when "0001011101111001" => data <= "001001";
        when "0001011101111010" => data <= "001001";
        when "0001011101111011" => data <= "001001";
        when "0001011101111100" => data <= "001001";
        when "0001011101111101" => data <= "001001";
        when "0001011101111110" => data <= "001001";
        when "0001011101111111" => data <= "001001";
        when "0001011110000000" => data <= "001001";
        when "0001011110000001" => data <= "001001";
        when "0001011110000010" => data <= "001001";
        when "0001011110000011" => data <= "110000";
        when "0001011110000100" => data <= "110000";
        when "0001011110001111" => data <= "111111";
        when "0001011110010011" => data <= "111111";
        when "0001011110010111" => data <= "111111";
        when "0001011110011110" => data <= "110000";
        when "0001011110011111" => data <= "110000";
        when "0001100000000000" => data <= "110000";
        when "0001100000000001" => data <= "110000";
        when "0001100000011001" => data <= "110000";
        when "0001100000011010" => data <= "110000";
        when "0001100000011011" => data <= "001001";
        when "0001100000011100" => data <= "001001";
        when "0001100000011101" => data <= "001001";
        when "0001100000011110" => data <= "001001";
        when "0001100000011111" => data <= "001001";
        when "0001100000100000" => data <= "001001";
        when "0001100000100001" => data <= "001001";
        when "0001100000100010" => data <= "001001";
        when "0001100000100011" => data <= "001001";
        when "0001100000100100" => data <= "001001";
        when "0001100000100101" => data <= "001001";
        when "0001100000100110" => data <= "001001";
        when "0001100000100111" => data <= "001001";
        when "0001100000101000" => data <= "001001";
        when "0001100000101001" => data <= "001001";
        when "0001100000101010" => data <= "001001";
        when "0001100000101011" => data <= "001001";
        when "0001100000101100" => data <= "001001";
        when "0001100000101101" => data <= "001001";
        when "0001100000101110" => data <= "001001";
        when "0001100000101111" => data <= "110000";
        when "0001100000110000" => data <= "110000";
        when "0001100001000101" => data <= "110000";
        when "0001100001000110" => data <= "110000";
        when "0001100001000111" => data <= "110000";
        when "0001100001001000" => data <= "110000";
        when "0001100001001001" => data <= "110000";
        when "0001100001010010" => data <= "110000";
        when "0001100001010011" => data <= "110000";
        when "0001100001010100" => data <= "110000";
        when "0001100001010101" => data <= "110000";
        when "0001100001010110" => data <= "110000";
        when "0001100001010111" => data <= "110000";
        when "0001100001110000" => data <= "110000";
        when "0001100001110001" => data <= "001001";
        when "0001100001110010" => data <= "001001";
        when "0001100001110011" => data <= "001001";
        when "0001100001110100" => data <= "001001";
        when "0001100001110101" => data <= "001001";
        when "0001100001110110" => data <= "001001";
        when "0001100001110111" => data <= "001001";
        when "0001100001111000" => data <= "001001";
        when "0001100001111001" => data <= "001001";
        when "0001100001111010" => data <= "001001";
        when "0001100001111011" => data <= "001001";
        when "0001100001111100" => data <= "001001";
        when "0001100001111101" => data <= "001001";
        when "0001100001111110" => data <= "001001";
        when "0001100001111111" => data <= "001001";
        when "0001100010000000" => data <= "001001";
        when "0001100010000001" => data <= "001001";
        when "0001100010000010" => data <= "001001";
        when "0001100010000011" => data <= "001001";
        when "0001100010000100" => data <= "001001";
        when "0001100010000101" => data <= "110000";
        when "0001100010000110" => data <= "110000";
        when "0001100010000111" => data <= "110000";
        when "0001100010011110" => data <= "110000";
        when "0001100010011111" => data <= "110000";
        when "0001100100000000" => data <= "110000";
        when "0001100100000001" => data <= "110000";
        when "0001100100010110" => data <= "110000";
        when "0001100100010111" => data <= "110000";
        when "0001100100011000" => data <= "110000";
        when "0001100100011001" => data <= "001001";
        when "0001100100011010" => data <= "001001";
        when "0001100100011011" => data <= "001001";
        when "0001100100011100" => data <= "001001";
        when "0001100100011101" => data <= "001001";
        when "0001100100011110" => data <= "001001";
        when "0001100100011111" => data <= "001001";
        when "0001100100100000" => data <= "001001";
        when "0001100100100001" => data <= "001001";
        when "0001100100100010" => data <= "001001";
        when "0001100100100011" => data <= "001001";
        when "0001100100100100" => data <= "001001";
        when "0001100100100101" => data <= "001001";
        when "0001100100100110" => data <= "001001";
        when "0001100100100111" => data <= "001001";
        when "0001100100101000" => data <= "001001";
        when "0001100100101001" => data <= "001001";
        when "0001100100101010" => data <= "001001";
        when "0001100100101011" => data <= "001001";
        when "0001100100101100" => data <= "001001";
        when "0001100100101101" => data <= "001001";
        when "0001100100101110" => data <= "110000";
        when "0001100101000101" => data <= "110000";
        when "0001100101000110" => data <= "110000";
        when "0001100101000111" => data <= "110000";
        when "0001100101001000" => data <= "110000";
        when "0001100101001001" => data <= "110000";
        when "0001100101010010" => data <= "110000";
        when "0001100101010011" => data <= "110000";
        when "0001100101010100" => data <= "110000";
        when "0001100101010101" => data <= "110000";
        when "0001100101010110" => data <= "110000";
        when "0001100101010111" => data <= "110000";
        when "0001100101110001" => data <= "110000";
        when "0001100101110010" => data <= "110000";
        when "0001100101110011" => data <= "001001";
        when "0001100101110100" => data <= "001001";
        when "0001100101110101" => data <= "001001";
        when "0001100101110110" => data <= "001001";
        when "0001100101110111" => data <= "001001";
        when "0001100101111000" => data <= "001001";
        when "0001100101111001" => data <= "001001";
        when "0001100101111010" => data <= "001001";
        when "0001100101111011" => data <= "001001";
        when "0001100101111100" => data <= "001001";
        when "0001100101111101" => data <= "001001";
        when "0001100101111110" => data <= "001001";
        when "0001100101111111" => data <= "001001";
        when "0001100110000000" => data <= "001001";
        when "0001100110000001" => data <= "001001";
        when "0001100110000010" => data <= "001001";
        when "0001100110000011" => data <= "001001";
        when "0001100110000100" => data <= "001001";
        when "0001100110000101" => data <= "001001";
        when "0001100110000110" => data <= "001001";
        when "0001100110000111" => data <= "001001";
        when "0001100110001000" => data <= "110000";
        when "0001100110001001" => data <= "110000";
        when "0001100110011110" => data <= "110000";
        when "0001100110011111" => data <= "110000";
        when "0001101000000000" => data <= "110000";
        when "0001101000000001" => data <= "110000";
        when "0001101000010100" => data <= "110000";
        when "0001101000010101" => data <= "110000";
        when "0001101000010110" => data <= "001001";
        when "0001101000010111" => data <= "001001";
        when "0001101000011000" => data <= "001001";
        when "0001101000011001" => data <= "001001";
        when "0001101000011010" => data <= "001001";
        when "0001101000011011" => data <= "001001";
        when "0001101000011100" => data <= "001001";
        when "0001101000011101" => data <= "001001";
        when "0001101000011110" => data <= "001001";
        when "0001101000011111" => data <= "001001";
        when "0001101000100000" => data <= "001001";
        when "0001101000100001" => data <= "001001";
        when "0001101000100010" => data <= "001001";
        when "0001101000100011" => data <= "001001";
        when "0001101000100100" => data <= "001001";
        when "0001101000100101" => data <= "001001";
        when "0001101000100110" => data <= "001001";
        when "0001101000100111" => data <= "001001";
        when "0001101000101000" => data <= "001001";
        when "0001101000101001" => data <= "001001";
        when "0001101000101010" => data <= "001001";
        when "0001101000101011" => data <= "001001";
        when "0001101000101100" => data <= "001001";
        when "0001101000101101" => data <= "110000";
        when "0001101001000101" => data <= "110000";
        when "0001101001000110" => data <= "110000";
        when "0001101001000111" => data <= "110000";
        when "0001101001001000" => data <= "110000";
        when "0001101001001001" => data <= "110000";
        when "0001101001010011" => data <= "110000";
        when "0001101001010100" => data <= "110000";
        when "0001101001010101" => data <= "110000";
        when "0001101001010110" => data <= "110000";
        when "0001101001110011" => data <= "110000";
        when "0001101001110100" => data <= "001001";
        when "0001101001110101" => data <= "001001";
        when "0001101001110110" => data <= "001001";
        when "0001101001110111" => data <= "001001";
        when "0001101001111000" => data <= "001001";
        when "0001101001111001" => data <= "001001";
        when "0001101001111010" => data <= "001001";
        when "0001101001111011" => data <= "001001";
        when "0001101001111100" => data <= "001001";
        when "0001101001111101" => data <= "001001";
        when "0001101001111110" => data <= "001001";
        when "0001101001111111" => data <= "001001";
        when "0001101010000000" => data <= "001001";
        when "0001101010000001" => data <= "001001";
        when "0001101010000010" => data <= "001001";
        when "0001101010000011" => data <= "001001";
        when "0001101010000100" => data <= "001001";
        when "0001101010000101" => data <= "001001";
        when "0001101010000110" => data <= "001001";
        when "0001101010000111" => data <= "001001";
        when "0001101010001000" => data <= "001001";
        when "0001101010001001" => data <= "001001";
        when "0001101010001010" => data <= "110000";
        when "0001101010001011" => data <= "110000";
        when "0001101010011110" => data <= "110000";
        when "0001101010011111" => data <= "110000";
        when "0001101100000000" => data <= "110000";
        when "0001101100000001" => data <= "110000";
        when "0001101100010010" => data <= "110000";
        when "0001101100010011" => data <= "110000";
        when "0001101100010100" => data <= "001001";
        when "0001101100010101" => data <= "001001";
        when "0001101100010110" => data <= "001001";
        when "0001101100010111" => data <= "001001";
        when "0001101100011000" => data <= "001001";
        when "0001101100011001" => data <= "001001";
        when "0001101100011010" => data <= "001001";
        when "0001101100011011" => data <= "001001";
        when "0001101100011100" => data <= "001001";
        when "0001101100011101" => data <= "001001";
        when "0001101100011110" => data <= "001001";
        when "0001101100011111" => data <= "001001";
        when "0001101100100000" => data <= "001001";
        when "0001101100100001" => data <= "001001";
        when "0001101100100010" => data <= "001001";
        when "0001101100100011" => data <= "001001";
        when "0001101100100100" => data <= "001001";
        when "0001101100100101" => data <= "001001";
        when "0001101100100110" => data <= "001001";
        when "0001101100100111" => data <= "001001";
        when "0001101100101000" => data <= "001001";
        when "0001101100101001" => data <= "001001";
        when "0001101100101010" => data <= "001001";
        when "0001101100101011" => data <= "110000";
        when "0001101100101100" => data <= "110000";
        when "0001101101000110" => data <= "110000";
        when "0001101101000111" => data <= "110000";
        when "0001101101001000" => data <= "110000";
        when "0001101101110100" => data <= "110000";
        when "0001101101110101" => data <= "001001";
        when "0001101101110110" => data <= "001001";
        when "0001101101110111" => data <= "001001";
        when "0001101101111000" => data <= "001001";
        when "0001101101111001" => data <= "001001";
        when "0001101101111010" => data <= "001001";
        when "0001101101111011" => data <= "001001";
        when "0001101101111100" => data <= "001001";
        when "0001101101111101" => data <= "001001";
        when "0001101101111110" => data <= "001001";
        when "0001101101111111" => data <= "001001";
        when "0001101110000000" => data <= "001001";
        when "0001101110000001" => data <= "001001";
        when "0001101110000010" => data <= "001001";
        when "0001101110000011" => data <= "001001";
        when "0001101110000100" => data <= "001001";
        when "0001101110000101" => data <= "001001";
        when "0001101110000110" => data <= "001001";
        when "0001101110000111" => data <= "001001";
        when "0001101110001000" => data <= "001001";
        when "0001101110001001" => data <= "001001";
        when "0001101110001010" => data <= "001001";
        when "0001101110001011" => data <= "001001";
        when "0001101110001100" => data <= "110000";
        when "0001101110001101" => data <= "110000";
        when "0001101110011110" => data <= "110000";
        when "0001101110011111" => data <= "110000";
        when "0001110000000000" => data <= "110000";
        when "0001110000000001" => data <= "110000";
        when "0001110000010000" => data <= "110000";
        when "0001110000010001" => data <= "110000";
        when "0001110000010010" => data <= "001001";
        when "0001110000010011" => data <= "001001";
        when "0001110000010100" => data <= "001001";
        when "0001110000010101" => data <= "001001";
        when "0001110000010110" => data <= "001001";
        when "0001110000010111" => data <= "001001";
        when "0001110000011000" => data <= "001001";
        when "0001110000011001" => data <= "001001";
        when "0001110000011010" => data <= "001001";
        when "0001110000011011" => data <= "001001";
        when "0001110000011100" => data <= "001001";
        when "0001110000011101" => data <= "001001";
        when "0001110000011110" => data <= "001001";
        when "0001110000011111" => data <= "001001";
        when "0001110000100000" => data <= "001001";
        when "0001110000100001" => data <= "001001";
        when "0001110000100010" => data <= "001001";
        when "0001110000100011" => data <= "001001";
        when "0001110000100100" => data <= "001001";
        when "0001110000100101" => data <= "001001";
        when "0001110000100110" => data <= "001001";
        when "0001110000100111" => data <= "001001";
        when "0001110000101000" => data <= "001001";
        when "0001110000101001" => data <= "001001";
        when "0001110000101010" => data <= "110000";
        when "0001110001110101" => data <= "110000";
        when "0001110001110110" => data <= "110000";
        when "0001110001110111" => data <= "001001";
        when "0001110001111000" => data <= "001001";
        when "0001110001111001" => data <= "001001";
        when "0001110001111010" => data <= "001001";
        when "0001110001111011" => data <= "001001";
        when "0001110001111100" => data <= "001001";
        when "0001110001111101" => data <= "001001";
        when "0001110001111110" => data <= "001001";
        when "0001110001111111" => data <= "001001";
        when "0001110010000000" => data <= "001001";
        when "0001110010000001" => data <= "001001";
        when "0001110010000010" => data <= "001001";
        when "0001110010000011" => data <= "001001";
        when "0001110010000100" => data <= "001001";
        when "0001110010000101" => data <= "001001";
        when "0001110010000110" => data <= "001001";
        when "0001110010000111" => data <= "001001";
        when "0001110010001000" => data <= "001001";
        when "0001110010001001" => data <= "001001";
        when "0001110010001010" => data <= "001001";
        when "0001110010001011" => data <= "001001";
        when "0001110010001100" => data <= "001001";
        when "0001110010001101" => data <= "001001";
        when "0001110010001110" => data <= "110000";
        when "0001110010001111" => data <= "110000";
        when "0001110010010000" => data <= "110000";
        when "0001110010011110" => data <= "110000";
        when "0001110010011111" => data <= "110000";
        when "0001110100000000" => data <= "110000";
        when "0001110100000001" => data <= "110000";
        when "0001110100001101" => data <= "110000";
        when "0001110100001110" => data <= "110000";
        when "0001110100001111" => data <= "110000";
        when "0001110100010000" => data <= "001001";
        when "0001110100010001" => data <= "001001";
        when "0001110100010010" => data <= "001001";
        when "0001110100010011" => data <= "001001";
        when "0001110100010100" => data <= "001001";
        when "0001110100010101" => data <= "001001";
        when "0001110100010110" => data <= "001001";
        when "0001110100010111" => data <= "001001";
        when "0001110100011000" => data <= "001001";
        when "0001110100011001" => data <= "001001";
        when "0001110100011010" => data <= "001001";
        when "0001110100011011" => data <= "001001";
        when "0001110100011100" => data <= "001001";
        when "0001110100011101" => data <= "001001";
        when "0001110100011110" => data <= "001001";
        when "0001110100011111" => data <= "001001";
        when "0001110100100000" => data <= "001001";
        when "0001110100100001" => data <= "001001";
        when "0001110100100010" => data <= "001001";
        when "0001110100100011" => data <= "001001";
        when "0001110100100100" => data <= "001001";
        when "0001110100100101" => data <= "001001";
        when "0001110100100110" => data <= "001001";
        when "0001110100100111" => data <= "001001";
        when "0001110100101000" => data <= "001001";
        when "0001110100101001" => data <= "110000";
        when "0001110101110111" => data <= "110000";
        when "0001110101111000" => data <= "001001";
        when "0001110101111001" => data <= "001001";
        when "0001110101111010" => data <= "001001";
        when "0001110101111011" => data <= "001001";
        when "0001110101111100" => data <= "001001";
        when "0001110101111101" => data <= "001001";
        when "0001110101111110" => data <= "001001";
        when "0001110101111111" => data <= "001001";
        when "0001110110000000" => data <= "001001";
        when "0001110110000001" => data <= "001001";
        when "0001110110000010" => data <= "001001";
        when "0001110110000011" => data <= "001001";
        when "0001110110000100" => data <= "001001";
        when "0001110110000101" => data <= "001001";
        when "0001110110000110" => data <= "001001";
        when "0001110110000111" => data <= "001001";
        when "0001110110001000" => data <= "001001";
        when "0001110110001001" => data <= "001001";
        when "0001110110001010" => data <= "001001";
        when "0001110110001011" => data <= "001001";
        when "0001110110001100" => data <= "001001";
        when "0001110110001101" => data <= "001001";
        when "0001110110001110" => data <= "001001";
        when "0001110110001111" => data <= "001001";
        when "0001110110010000" => data <= "001001";
        when "0001110110010001" => data <= "110000";
        when "0001110110010010" => data <= "110000";
        when "0001110110011110" => data <= "110000";
        when "0001110110011111" => data <= "110000";
        when "0001111000000000" => data <= "110000";
        when "0001111000000001" => data <= "110000";
        when "0001111000001011" => data <= "110000";
        when "0001111000001100" => data <= "110000";
        when "0001111000001101" => data <= "001001";
        when "0001111000001110" => data <= "001001";
        when "0001111000001111" => data <= "001001";
        when "0001111000010000" => data <= "001001";
        when "0001111000010001" => data <= "001001";
        when "0001111000010010" => data <= "001001";
        when "0001111000010011" => data <= "001001";
        when "0001111000010100" => data <= "001001";
        when "0001111000010101" => data <= "001001";
        when "0001111000010110" => data <= "001001";
        when "0001111000010111" => data <= "001001";
        when "0001111000011000" => data <= "001001";
        when "0001111000011001" => data <= "001001";
        when "0001111000011010" => data <= "001001";
        when "0001111000011011" => data <= "001001";
        when "0001111000011100" => data <= "001001";
        when "0001111000011101" => data <= "001001";
        when "0001111000011110" => data <= "001001";
        when "0001111000011111" => data <= "001001";
        when "0001111000100000" => data <= "001001";
        when "0001111000100001" => data <= "001001";
        when "0001111000100010" => data <= "001001";
        when "0001111000100011" => data <= "001001";
        when "0001111000100100" => data <= "001001";
        when "0001111000100101" => data <= "001001";
        when "0001111000100110" => data <= "001001";
        when "0001111000100111" => data <= "110000";
        when "0001111000101000" => data <= "110000";
        when "0001111001111000" => data <= "110000";
        when "0001111001111001" => data <= "001001";
        when "0001111001111010" => data <= "001001";
        when "0001111001111011" => data <= "001001";
        when "0001111001111100" => data <= "001001";
        when "0001111001111101" => data <= "001001";
        when "0001111001111110" => data <= "001001";
        when "0001111001111111" => data <= "001001";
        when "0001111010000000" => data <= "001001";
        when "0001111010000001" => data <= "001001";
        when "0001111010000010" => data <= "001001";
        when "0001111010000011" => data <= "001001";
        when "0001111010000100" => data <= "001001";
        when "0001111010000101" => data <= "001001";
        when "0001111010000110" => data <= "001001";
        when "0001111010000111" => data <= "001001";
        when "0001111010001000" => data <= "001001";
        when "0001111010001001" => data <= "001001";
        when "0001111010001010" => data <= "001001";
        when "0001111010001011" => data <= "001001";
        when "0001111010001100" => data <= "001001";
        when "0001111010001101" => data <= "001001";
        when "0001111010001110" => data <= "001001";
        when "0001111010001111" => data <= "001001";
        when "0001111010010000" => data <= "001001";
        when "0001111010010001" => data <= "001001";
        when "0001111010010010" => data <= "001001";
        when "0001111010010011" => data <= "110000";
        when "0001111010010100" => data <= "110000";
        when "0001111010011110" => data <= "110000";
        when "0001111010011111" => data <= "110000";
        when "0001111100000000" => data <= "110000";
        when "0001111100000001" => data <= "110000";
        when "0001111100001011" => data <= "110000";
        when "0001111100001100" => data <= "001001";
        when "0001111100001101" => data <= "001001";
        when "0001111100001110" => data <= "001001";
        when "0001111100001111" => data <= "001001";
        when "0001111100010000" => data <= "001001";
        when "0001111100010001" => data <= "001001";
        when "0001111100010010" => data <= "001001";
        when "0001111100010011" => data <= "001001";
        when "0001111100010100" => data <= "001001";
        when "0001111100010101" => data <= "001001";
        when "0001111100010110" => data <= "001001";
        when "0001111100010111" => data <= "001001";
        when "0001111100011000" => data <= "001001";
        when "0001111100011001" => data <= "001001";
        when "0001111100011010" => data <= "001001";
        when "0001111100011011" => data <= "001001";
        when "0001111100011100" => data <= "001001";
        when "0001111100011101" => data <= "001001";
        when "0001111100011110" => data <= "001001";
        when "0001111100011111" => data <= "001001";
        when "0001111100100000" => data <= "001001";
        when "0001111100100001" => data <= "001001";
        when "0001111100100010" => data <= "001001";
        when "0001111100100011" => data <= "001001";
        when "0001111100100100" => data <= "001001";
        when "0001111100100101" => data <= "001001";
        when "0001111100100110" => data <= "110000";
        when "0001111101111001" => data <= "110000";
        when "0001111101111010" => data <= "110000";
        when "0001111101111011" => data <= "001001";
        when "0001111101111100" => data <= "001001";
        when "0001111101111101" => data <= "001001";
        when "0001111101111110" => data <= "001001";
        when "0001111101111111" => data <= "001001";
        when "0001111110000000" => data <= "001001";
        when "0001111110000001" => data <= "001001";
        when "0001111110000010" => data <= "001001";
        when "0001111110000011" => data <= "001001";
        when "0001111110000100" => data <= "001001";
        when "0001111110000101" => data <= "001001";
        when "0001111110000110" => data <= "001001";
        when "0001111110000111" => data <= "001001";
        when "0001111110001000" => data <= "001001";
        when "0001111110001001" => data <= "001001";
        when "0001111110001010" => data <= "001001";
        when "0001111110001011" => data <= "001001";
        when "0001111110001100" => data <= "001001";
        when "0001111110001101" => data <= "001001";
        when "0001111110001110" => data <= "001001";
        when "0001111110001111" => data <= "001001";
        when "0001111110010000" => data <= "001001";
        when "0001111110010001" => data <= "001001";
        when "0001111110010010" => data <= "001001";
        when "0001111110010011" => data <= "001001";
        when "0001111110010100" => data <= "110000";
        when "0001111110011110" => data <= "110000";
        when "0001111110011111" => data <= "110000";
        when "0010000000000000" => data <= "110000";
        when "0010000000000001" => data <= "110000";
        when "0010000000001011" => data <= "110000";
        when "0010000000001100" => data <= "001001";
        when "0010000000001101" => data <= "001001";
        when "0010000000001110" => data <= "001001";
        when "0010000000001111" => data <= "001001";
        when "0010000000010000" => data <= "001001";
        when "0010000000010001" => data <= "001001";
        when "0010000000010010" => data <= "001001";
        when "0010000000010011" => data <= "001001";
        when "0010000000010100" => data <= "001001";
        when "0010000000010101" => data <= "001001";
        when "0010000000010110" => data <= "001001";
        when "0010000000010111" => data <= "001001";
        when "0010000000011000" => data <= "001001";
        when "0010000000011001" => data <= "001001";
        when "0010000000011010" => data <= "001001";
        when "0010000000011011" => data <= "001001";
        when "0010000000011100" => data <= "001001";
        when "0010000000011101" => data <= "001001";
        when "0010000000011110" => data <= "001001";
        when "0010000000011111" => data <= "001001";
        when "0010000000100000" => data <= "001001";
        when "0010000000100001" => data <= "001001";
        when "0010000000100010" => data <= "001001";
        when "0010000000100011" => data <= "001001";
        when "0010000000100100" => data <= "110000";
        when "0010000000100101" => data <= "110000";
        when "0010000001111011" => data <= "110000";
        when "0010000001111100" => data <= "001001";
        when "0010000001111101" => data <= "001001";
        when "0010000001111110" => data <= "001001";
        when "0010000001111111" => data <= "001001";
        when "0010000010000000" => data <= "001001";
        when "0010000010000001" => data <= "001001";
        when "0010000010000010" => data <= "001001";
        when "0010000010000011" => data <= "001001";
        when "0010000010000100" => data <= "001001";
        when "0010000010000101" => data <= "001001";
        when "0010000010000110" => data <= "001001";
        when "0010000010000111" => data <= "001001";
        when "0010000010001000" => data <= "001001";
        when "0010000010001001" => data <= "001001";
        when "0010000010001010" => data <= "001001";
        when "0010000010001011" => data <= "001001";
        when "0010000010001100" => data <= "001001";
        when "0010000010001101" => data <= "001001";
        when "0010000010001110" => data <= "001001";
        when "0010000010001111" => data <= "001001";
        when "0010000010010000" => data <= "001001";
        when "0010000010010001" => data <= "001001";
        when "0010000010010010" => data <= "001001";
        when "0010000010010011" => data <= "001001";
        when "0010000010010100" => data <= "110000";
        when "0010000010011110" => data <= "110000";
        when "0010000010011111" => data <= "110000";
        when "0010000100000000" => data <= "110000";
        when "0010000100000001" => data <= "110000";
        when "0010000100001011" => data <= "110000";
        when "0010000100001100" => data <= "001001";
        when "0010000100001101" => data <= "001001";
        when "0010000100001110" => data <= "001001";
        when "0010000100001111" => data <= "001001";
        when "0010000100010000" => data <= "001001";
        when "0010000100010001" => data <= "001001";
        when "0010000100010010" => data <= "001001";
        when "0010000100010011" => data <= "001001";
        when "0010000100010100" => data <= "001001";
        when "0010000100010101" => data <= "001001";
        when "0010000100010110" => data <= "001001";
        when "0010000100010111" => data <= "001001";
        when "0010000100011000" => data <= "001001";
        when "0010000100011001" => data <= "001001";
        when "0010000100011010" => data <= "001001";
        when "0010000100011011" => data <= "001001";
        when "0010000100011100" => data <= "001001";
        when "0010000100011101" => data <= "001001";
        when "0010000100011110" => data <= "001001";
        when "0010000100011111" => data <= "001001";
        when "0010000100100000" => data <= "001001";
        when "0010000100100001" => data <= "001001";
        when "0010000100100010" => data <= "001001";
        when "0010000100100011" => data <= "110000";
        when "0010000101111100" => data <= "110000";
        when "0010000101111101" => data <= "001001";
        when "0010000101111110" => data <= "001001";
        when "0010000101111111" => data <= "001001";
        when "0010000110000000" => data <= "001001";
        when "0010000110000001" => data <= "001001";
        when "0010000110000010" => data <= "001001";
        when "0010000110000011" => data <= "001001";
        when "0010000110000100" => data <= "001001";
        when "0010000110000101" => data <= "001001";
        when "0010000110000110" => data <= "001001";
        when "0010000110000111" => data <= "001001";
        when "0010000110001000" => data <= "001001";
        when "0010000110001001" => data <= "001001";
        when "0010000110001010" => data <= "001001";
        when "0010000110001011" => data <= "001001";
        when "0010000110001100" => data <= "001001";
        when "0010000110001101" => data <= "001001";
        when "0010000110001110" => data <= "001001";
        when "0010000110001111" => data <= "001001";
        when "0010000110010000" => data <= "001001";
        when "0010000110010001" => data <= "001001";
        when "0010000110010010" => data <= "001001";
        when "0010000110010011" => data <= "001001";
        when "0010000110010100" => data <= "110000";
        when "0010000110011110" => data <= "110000";
        when "0010000110011111" => data <= "110000";
        when "0010001000000000" => data <= "110000";
        when "0010001000000001" => data <= "110000";
        when "0010001000001011" => data <= "110000";
        when "0010001000001100" => data <= "001001";
        when "0010001000001101" => data <= "001001";
        when "0010001000001110" => data <= "001001";
        when "0010001000001111" => data <= "001001";
        when "0010001000010000" => data <= "001001";
        when "0010001000010001" => data <= "001001";
        when "0010001000010010" => data <= "001001";
        when "0010001000010011" => data <= "001001";
        when "0010001000010100" => data <= "001001";
        when "0010001000010101" => data <= "001001";
        when "0010001000010110" => data <= "001001";
        when "0010001000010111" => data <= "001001";
        when "0010001000011000" => data <= "001001";
        when "0010001000011001" => data <= "001001";
        when "0010001000011010" => data <= "001001";
        when "0010001000011011" => data <= "001001";
        when "0010001000011100" => data <= "001001";
        when "0010001000011101" => data <= "001001";
        when "0010001000011110" => data <= "001001";
        when "0010001000011111" => data <= "001001";
        when "0010001000100000" => data <= "001001";
        when "0010001000100001" => data <= "001001";
        when "0010001000100010" => data <= "110000";
        when "0010001001111101" => data <= "110000";
        when "0010001001111110" => data <= "110000";
        when "0010001001111111" => data <= "001001";
        when "0010001010000000" => data <= "001001";
        when "0010001010000001" => data <= "001001";
        when "0010001010000010" => data <= "001001";
        when "0010001010000011" => data <= "001001";
        when "0010001010000100" => data <= "001001";
        when "0010001010000101" => data <= "001001";
        when "0010001010000110" => data <= "001001";
        when "0010001010000111" => data <= "001001";
        when "0010001010001000" => data <= "001001";
        when "0010001010001001" => data <= "001001";
        when "0010001010001010" => data <= "001001";
        when "0010001010001011" => data <= "001001";
        when "0010001010001100" => data <= "001001";
        when "0010001010001101" => data <= "001001";
        when "0010001010001110" => data <= "001001";
        when "0010001010001111" => data <= "001001";
        when "0010001010010000" => data <= "001001";
        when "0010001010010001" => data <= "001001";
        when "0010001010010010" => data <= "001001";
        when "0010001010010011" => data <= "001001";
        when "0010001010010100" => data <= "110000";
        when "0010001010011110" => data <= "110000";
        when "0010001010011111" => data <= "110000";
        when "0010001100000000" => data <= "110000";
        when "0010001100000001" => data <= "110000";
        when "0010001100001011" => data <= "110000";
        when "0010001100001100" => data <= "001001";
        when "0010001100001101" => data <= "001001";
        when "0010001100001110" => data <= "001001";
        when "0010001100001111" => data <= "001001";
        when "0010001100010000" => data <= "001001";
        when "0010001100010001" => data <= "001001";
        when "0010001100010010" => data <= "001001";
        when "0010001100010011" => data <= "001001";
        when "0010001100010100" => data <= "001001";
        when "0010001100010101" => data <= "001001";
        when "0010001100010110" => data <= "001001";
        when "0010001100010111" => data <= "001001";
        when "0010001100011000" => data <= "001001";
        when "0010001100011001" => data <= "001001";
        when "0010001100011010" => data <= "001001";
        when "0010001100011011" => data <= "001001";
        when "0010001100011100" => data <= "001001";
        when "0010001100011101" => data <= "001001";
        when "0010001100011110" => data <= "001001";
        when "0010001100011111" => data <= "001001";
        when "0010001100100000" => data <= "110000";
        when "0010001100100001" => data <= "110000";
        when "0010001101111111" => data <= "110000";
        when "0010001110000000" => data <= "001001";
        when "0010001110000001" => data <= "001001";
        when "0010001110000010" => data <= "001001";
        when "0010001110000011" => data <= "001001";
        when "0010001110000100" => data <= "001001";
        when "0010001110000101" => data <= "001001";
        when "0010001110000110" => data <= "001001";
        when "0010001110000111" => data <= "001001";
        when "0010001110001000" => data <= "001001";
        when "0010001110001001" => data <= "001001";
        when "0010001110001010" => data <= "001001";
        when "0010001110001011" => data <= "001001";
        when "0010001110001100" => data <= "001001";
        when "0010001110001101" => data <= "001001";
        when "0010001110001110" => data <= "001001";
        when "0010001110001111" => data <= "001001";
        when "0010001110010000" => data <= "001001";
        when "0010001110010001" => data <= "001001";
        when "0010001110010010" => data <= "001001";
        when "0010001110010011" => data <= "001001";
        when "0010001110010100" => data <= "110000";
        when "0010001110011110" => data <= "110000";
        when "0010001110011111" => data <= "110000";
        when "0010010000000000" => data <= "110000";
        when "0010010000000001" => data <= "110000";
        when "0010010000001011" => data <= "110000";
        when "0010010000001100" => data <= "001001";
        when "0010010000001101" => data <= "001001";
        when "0010010000001110" => data <= "001001";
        when "0010010000001111" => data <= "001001";
        when "0010010000010000" => data <= "001001";
        when "0010010000010001" => data <= "001001";
        when "0010010000010010" => data <= "001001";
        when "0010010000010011" => data <= "001001";
        when "0010010000010100" => data <= "001001";
        when "0010010000010101" => data <= "001001";
        when "0010010000010110" => data <= "001001";
        when "0010010000010111" => data <= "001001";
        when "0010010000011000" => data <= "001001";
        when "0010010000011001" => data <= "001001";
        when "0010010000011010" => data <= "001001";
        when "0010010000011011" => data <= "001001";
        when "0010010000011100" => data <= "001001";
        when "0010010000011101" => data <= "001001";
        when "0010010000011110" => data <= "001001";
        when "0010010000011111" => data <= "110000";
        when "0010010010000000" => data <= "110000";
        when "0010010010000001" => data <= "001001";
        when "0010010010000010" => data <= "001001";
        when "0010010010000011" => data <= "001001";
        when "0010010010000100" => data <= "001001";
        when "0010010010000101" => data <= "001001";
        when "0010010010000110" => data <= "001001";
        when "0010010010000111" => data <= "001001";
        when "0010010010001000" => data <= "001001";
        when "0010010010001001" => data <= "001001";
        when "0010010010001010" => data <= "001001";
        when "0010010010001011" => data <= "001001";
        when "0010010010001100" => data <= "001001";
        when "0010010010001101" => data <= "001001";
        when "0010010010001110" => data <= "001001";
        when "0010010010001111" => data <= "001001";
        when "0010010010010000" => data <= "001001";
        when "0010010010010001" => data <= "001001";
        when "0010010010010010" => data <= "001001";
        when "0010010010010011" => data <= "001001";
        when "0010010010010100" => data <= "110000";
        when "0010010010011110" => data <= "110000";
        when "0010010010011111" => data <= "110000";
        when "0010010100000000" => data <= "110000";
        when "0010010100000001" => data <= "110000";
        when "0010010100001011" => data <= "110000";
        when "0010010100001100" => data <= "001001";
        when "0010010100001101" => data <= "001001";
        when "0010010100001110" => data <= "001001";
        when "0010010100001111" => data <= "001001";
        when "0010010100010000" => data <= "001001";
        when "0010010100010001" => data <= "001001";
        when "0010010100010010" => data <= "001001";
        when "0010010100010011" => data <= "001001";
        when "0010010100010100" => data <= "001001";
        when "0010010100010101" => data <= "001001";
        when "0010010100010110" => data <= "001001";
        when "0010010100010111" => data <= "001001";
        when "0010010100011000" => data <= "001001";
        when "0010010100011001" => data <= "001001";
        when "0010010100011010" => data <= "001001";
        when "0010010100011011" => data <= "001001";
        when "0010010100011100" => data <= "001001";
        when "0010010100011101" => data <= "001001";
        when "0010010100011110" => data <= "110000";
        when "0010010110000001" => data <= "110000";
        when "0010010110000010" => data <= "110000";
        when "0010010110000011" => data <= "001001";
        when "0010010110000100" => data <= "001001";
        when "0010010110000101" => data <= "001001";
        when "0010010110000110" => data <= "001001";
        when "0010010110000111" => data <= "001001";
        when "0010010110001000" => data <= "001001";
        when "0010010110001001" => data <= "001001";
        when "0010010110001010" => data <= "001001";
        when "0010010110001011" => data <= "001001";
        when "0010010110001100" => data <= "001001";
        when "0010010110001101" => data <= "001001";
        when "0010010110001110" => data <= "001001";
        when "0010010110001111" => data <= "001001";
        when "0010010110010000" => data <= "001001";
        when "0010010110010001" => data <= "001001";
        when "0010010110010010" => data <= "001001";
        when "0010010110010011" => data <= "001001";
        when "0010010110010100" => data <= "110000";
        when "0010010110011110" => data <= "110000";
        when "0010010110011111" => data <= "110000";
        when "0010011000000000" => data <= "110000";
        when "0010011000000001" => data <= "110000";
        when "0010011000001011" => data <= "110000";
        when "0010011000001100" => data <= "001001";
        when "0010011000001101" => data <= "001001";
        when "0010011000001110" => data <= "001001";
        when "0010011000001111" => data <= "001001";
        when "0010011000010000" => data <= "001001";
        when "0010011000010001" => data <= "001001";
        when "0010011000010010" => data <= "001001";
        when "0010011000010011" => data <= "001001";
        when "0010011000010100" => data <= "001001";
        when "0010011000010101" => data <= "001001";
        when "0010011000010110" => data <= "001001";
        when "0010011000010111" => data <= "001001";
        when "0010011000011000" => data <= "001001";
        when "0010011000011001" => data <= "001001";
        when "0010011000011010" => data <= "001001";
        when "0010011000011011" => data <= "001001";
        when "0010011000011100" => data <= "110000";
        when "0010011000011101" => data <= "110000";
        when "0010011010000011" => data <= "110000";
        when "0010011010000100" => data <= "001001";
        when "0010011010000101" => data <= "001001";
        when "0010011010000110" => data <= "001001";
        when "0010011010000111" => data <= "001001";
        when "0010011010001000" => data <= "001001";
        when "0010011010001001" => data <= "001001";
        when "0010011010001010" => data <= "001001";
        when "0010011010001011" => data <= "001001";
        when "0010011010001100" => data <= "001001";
        when "0010011010001101" => data <= "001001";
        when "0010011010001110" => data <= "001001";
        when "0010011010001111" => data <= "001001";
        when "0010011010010000" => data <= "001001";
        when "0010011010010001" => data <= "001001";
        when "0010011010010010" => data <= "001001";
        when "0010011010010011" => data <= "001001";
        when "0010011010010100" => data <= "110000";
        when "0010011010011110" => data <= "110000";
        when "0010011010011111" => data <= "110000";
        when "0010011100000000" => data <= "110000";
        when "0010011100000001" => data <= "110000";
        when "0010011100001011" => data <= "110000";
        when "0010011100001100" => data <= "001001";
        when "0010011100001101" => data <= "001001";
        when "0010011100001110" => data <= "001001";
        when "0010011100001111" => data <= "001001";
        when "0010011100010000" => data <= "001001";
        when "0010011100010001" => data <= "001001";
        when "0010011100010010" => data <= "001001";
        when "0010011100010011" => data <= "001001";
        when "0010011100010100" => data <= "001001";
        when "0010011100010101" => data <= "001001";
        when "0010011100010110" => data <= "001001";
        when "0010011100010111" => data <= "001001";
        when "0010011100011000" => data <= "001001";
        when "0010011100011001" => data <= "001001";
        when "0010011100011010" => data <= "001001";
        when "0010011100011011" => data <= "110000";
        when "0010011110000100" => data <= "110000";
        when "0010011110000101" => data <= "001001";
        when "0010011110000110" => data <= "001001";
        when "0010011110000111" => data <= "001001";
        when "0010011110001000" => data <= "001001";
        when "0010011110001001" => data <= "001001";
        when "0010011110001010" => data <= "001001";
        when "0010011110001011" => data <= "001001";
        when "0010011110001100" => data <= "001001";
        when "0010011110001101" => data <= "001001";
        when "0010011110001110" => data <= "001001";
        when "0010011110001111" => data <= "001001";
        when "0010011110010000" => data <= "001001";
        when "0010011110010001" => data <= "001001";
        when "0010011110010010" => data <= "001001";
        when "0010011110010011" => data <= "001001";
        when "0010011110010100" => data <= "110000";
        when "0010011110011110" => data <= "110000";
        when "0010011110011111" => data <= "110000";
        when "0010100000000000" => data <= "110000";
        when "0010100000000001" => data <= "110000";
        when "0010100000001011" => data <= "110000";
        when "0010100000001100" => data <= "001001";
        when "0010100000001101" => data <= "001001";
        when "0010100000001110" => data <= "001001";
        when "0010100000001111" => data <= "001001";
        when "0010100000010000" => data <= "001001";
        when "0010100000010001" => data <= "001001";
        when "0010100000010010" => data <= "001001";
        when "0010100000010011" => data <= "001001";
        when "0010100000010100" => data <= "001001";
        when "0010100000010101" => data <= "001001";
        when "0010100000010110" => data <= "001001";
        when "0010100000010111" => data <= "001001";
        when "0010100000011000" => data <= "001001";
        when "0010100000011001" => data <= "001001";
        when "0010100000011010" => data <= "110000";
        when "0010100000011111" => data <= "110000";
        when "0010100000100101" => data <= "110000";
        when "0010100001001111" => data <= "110000";
        when "0010100001010101" => data <= "110000";
        when "0010100001100001" => data <= "110000";
        when "0010100010000101" => data <= "110000";
        when "0010100010000110" => data <= "110000";
        when "0010100010000111" => data <= "001001";
        when "0010100010001000" => data <= "001001";
        when "0010100010001001" => data <= "001001";
        when "0010100010001010" => data <= "001001";
        when "0010100010001011" => data <= "001001";
        when "0010100010001100" => data <= "001001";
        when "0010100010001101" => data <= "001001";
        when "0010100010001110" => data <= "001001";
        when "0010100010001111" => data <= "001001";
        when "0010100010010000" => data <= "001001";
        when "0010100010010001" => data <= "001001";
        when "0010100010010010" => data <= "001001";
        when "0010100010010011" => data <= "001001";
        when "0010100010010100" => data <= "110000";
        when "0010100010011110" => data <= "110000";
        when "0010100010011111" => data <= "110000";
        when "0010100100000000" => data <= "110000";
        when "0010100100000001" => data <= "110000";
        when "0010100100001011" => data <= "110000";
        when "0010100100001100" => data <= "001001";
        when "0010100100001101" => data <= "001001";
        when "0010100100001110" => data <= "001001";
        when "0010100100001111" => data <= "001001";
        when "0010100100010000" => data <= "001001";
        when "0010100100010001" => data <= "001001";
        when "0010100100010010" => data <= "001001";
        when "0010100100010011" => data <= "001001";
        when "0010100100010100" => data <= "001001";
        when "0010100100010101" => data <= "001001";
        when "0010100100010110" => data <= "001001";
        when "0010100100010111" => data <= "001001";
        when "0010100100011000" => data <= "110000";
        when "0010100100011001" => data <= "110000";
        when "0010100100011110" => data <= "110000";
        when "0010100100011111" => data <= "110000";
        when "0010100100100100" => data <= "110000";
        when "0010100100100101" => data <= "110000";
        when "0010100100101111" => data <= "110000";
        when "0010100100110000" => data <= "110000";
        when "0010100100111011" => data <= "110000";
        when "0010100100111100" => data <= "110000";
        when "0010100101001110" => data <= "110000";
        when "0010100101001111" => data <= "110000";
        when "0010100101010100" => data <= "110000";
        when "0010100101010101" => data <= "110000";
        when "0010100101100000" => data <= "110000";
        when "0010100101100001" => data <= "110000";
        when "0010100101100101" => data <= "110000";
        when "0010100101100110" => data <= "110000";
        when "0010100110000111" => data <= "110000";
        when "0010100110001000" => data <= "001001";
        when "0010100110001001" => data <= "001001";
        when "0010100110001010" => data <= "001001";
        when "0010100110001011" => data <= "001001";
        when "0010100110001100" => data <= "001001";
        when "0010100110001101" => data <= "001001";
        when "0010100110001110" => data <= "001001";
        when "0010100110001111" => data <= "001001";
        when "0010100110010000" => data <= "001001";
        when "0010100110010001" => data <= "001001";
        when "0010100110010010" => data <= "001001";
        when "0010100110010011" => data <= "001001";
        when "0010100110010100" => data <= "110000";
        when "0010100110011110" => data <= "110000";
        when "0010100110011111" => data <= "110000";
        when "0010101000000000" => data <= "110000";
        when "0010101000000001" => data <= "110000";
        when "0010101000001011" => data <= "110000";
        when "0010101000001100" => data <= "001001";
        when "0010101000001101" => data <= "001001";
        when "0010101000001110" => data <= "001001";
        when "0010101000001111" => data <= "001001";
        when "0010101000010000" => data <= "001001";
        when "0010101000010001" => data <= "001001";
        when "0010101000010010" => data <= "001001";
        when "0010101000010011" => data <= "001001";
        when "0010101000010100" => data <= "001001";
        when "0010101000010101" => data <= "001001";
        when "0010101000010110" => data <= "001001";
        when "0010101000010111" => data <= "110000";
        when "0010101000011110" => data <= "110000";
        when "0010101000011111" => data <= "110000";
        when "0010101000100100" => data <= "110000";
        when "0010101000100101" => data <= "110000";
        when "0010101000101111" => data <= "110000";
        when "0010101000110000" => data <= "110000";
        when "0010101000111011" => data <= "110000";
        when "0010101000111100" => data <= "110000";
        when "0010101001001110" => data <= "110000";
        when "0010101001001111" => data <= "110000";
        when "0010101001010100" => data <= "110000";
        when "0010101001010101" => data <= "110000";
        when "0010101001100000" => data <= "110000";
        when "0010101001100001" => data <= "110000";
        when "0010101001100101" => data <= "110000";
        when "0010101001100110" => data <= "110000";
        when "0010101010001000" => data <= "110000";
        when "0010101010001001" => data <= "001001";
        when "0010101010001010" => data <= "001001";
        when "0010101010001011" => data <= "001001";
        when "0010101010001100" => data <= "001001";
        when "0010101010001101" => data <= "001001";
        when "0010101010001110" => data <= "001001";
        when "0010101010001111" => data <= "001001";
        when "0010101010010000" => data <= "001001";
        when "0010101010010001" => data <= "001001";
        when "0010101010010010" => data <= "001001";
        when "0010101010010011" => data <= "001001";
        when "0010101010010100" => data <= "110000";
        when "0010101010011110" => data <= "110000";
        when "0010101010011111" => data <= "110000";
        when "0010101100000000" => data <= "110000";
        when "0010101100000001" => data <= "110000";
        when "0010101100001011" => data <= "110000";
        when "0010101100001100" => data <= "001001";
        when "0010101100001101" => data <= "001001";
        when "0010101100001110" => data <= "001001";
        when "0010101100001111" => data <= "001001";
        when "0010101100010000" => data <= "001001";
        when "0010101100010001" => data <= "001001";
        when "0010101100010010" => data <= "001001";
        when "0010101100010011" => data <= "001001";
        when "0010101100010100" => data <= "001001";
        when "0010101100010101" => data <= "001001";
        when "0010101100010110" => data <= "110000";
        when "0010101100011110" => data <= "110000";
        when "0010101100011111" => data <= "110000";
        when "0010101100100100" => data <= "110000";
        when "0010101100100101" => data <= "110000";
        when "0010101100101111" => data <= "110000";
        when "0010101100110000" => data <= "110000";
        when "0010101100111011" => data <= "110000";
        when "0010101100111100" => data <= "110000";
        when "0010101101001110" => data <= "110000";
        when "0010101101001111" => data <= "110000";
        when "0010101101010100" => data <= "110000";
        when "0010101101010101" => data <= "110000";
        when "0010101101100000" => data <= "110000";
        when "0010101101100001" => data <= "110000";
        when "0010101101100110" => data <= "110000";
        when "0010101101101010" => data <= "110000";
        when "0010101101101011" => data <= "110000";
        when "0010101110001001" => data <= "110000";
        when "0010101110001010" => data <= "110000";
        when "0010101110001011" => data <= "001001";
        when "0010101110001100" => data <= "001001";
        when "0010101110001101" => data <= "001001";
        when "0010101110001110" => data <= "001001";
        when "0010101110001111" => data <= "001001";
        when "0010101110010000" => data <= "001001";
        when "0010101110010001" => data <= "001001";
        when "0010101110010010" => data <= "001001";
        when "0010101110010011" => data <= "001001";
        when "0010101110010100" => data <= "110000";
        when "0010101110011110" => data <= "110000";
        when "0010101110011111" => data <= "110000";
        when "0010110000000000" => data <= "110000";
        when "0010110000000001" => data <= "110000";
        when "0010110000001011" => data <= "110000";
        when "0010110000001100" => data <= "001001";
        when "0010110000001101" => data <= "001001";
        when "0010110000001110" => data <= "001001";
        when "0010110000001111" => data <= "001001";
        when "0010110000010000" => data <= "001001";
        when "0010110000010001" => data <= "001001";
        when "0010110000010010" => data <= "001001";
        when "0010110000010011" => data <= "001001";
        when "0010110000010100" => data <= "110000";
        when "0010110000010101" => data <= "110000";
        when "0010110000011110" => data <= "110000";
        when "0010110000011111" => data <= "110000";
        when "0010110000100000" => data <= "110000";
        when "0010110000100100" => data <= "110000";
        when "0010110000100101" => data <= "110000";
        when "0010110000110000" => data <= "110000";
        when "0010110000110100" => data <= "110000";
        when "0010110000111011" => data <= "110000";
        when "0010110001001110" => data <= "110000";
        when "0010110001001111" => data <= "110000";
        when "0010110001010000" => data <= "110000";
        when "0010110001010100" => data <= "110000";
        when "0010110001010101" => data <= "110000";
        when "0010110001011111" => data <= "110000";
        when "0010110001100000" => data <= "110000";
        when "0010110001100001" => data <= "110000";
        when "0010110001100010" => data <= "110000";
        when "0010110001100011" => data <= "110000";
        when "0010110001100110" => data <= "110000";
        when "0010110001101001" => data <= "110000";
        when "0010110001101010" => data <= "110000";
        when "0010110010001011" => data <= "110000";
        when "0010110010001100" => data <= "001001";
        when "0010110010001101" => data <= "001001";
        when "0010110010001110" => data <= "001001";
        when "0010110010001111" => data <= "001001";
        when "0010110010010000" => data <= "001001";
        when "0010110010010001" => data <= "001001";
        when "0010110010010010" => data <= "001001";
        when "0010110010010011" => data <= "001001";
        when "0010110010010100" => data <= "110000";
        when "0010110010011110" => data <= "110000";
        when "0010110010011111" => data <= "110000";
        when "0010110100000000" => data <= "110000";
        when "0010110100000001" => data <= "110000";
        when "0010110100001011" => data <= "110000";
        when "0010110100001100" => data <= "001001";
        when "0010110100001101" => data <= "001001";
        when "0010110100001110" => data <= "001001";
        when "0010110100001111" => data <= "001001";
        when "0010110100010000" => data <= "001001";
        when "0010110100010001" => data <= "001001";
        when "0010110100010010" => data <= "001001";
        when "0010110100010011" => data <= "110000";
        when "0010110100011110" => data <= "110000";
        when "0010110100011111" => data <= "110000";
        when "0010110100100000" => data <= "110000";
        when "0010110100100001" => data <= "110000";
        when "0010110100100010" => data <= "110000";
        when "0010110100100011" => data <= "110000";
        when "0010110100100100" => data <= "110000";
        when "0010110100100101" => data <= "110000";
        when "0010110100110000" => data <= "110000";
        when "0010110100110011" => data <= "110000";
        when "0010110100110100" => data <= "110000";
        when "0010110100111011" => data <= "110000";
        when "0010110101001110" => data <= "110000";
        when "0010110101001111" => data <= "110000";
        when "0010110101010000" => data <= "110000";
        when "0010110101010001" => data <= "110000";
        when "0010110101010010" => data <= "110000";
        when "0010110101010011" => data <= "110000";
        when "0010110101010100" => data <= "110000";
        when "0010110101010101" => data <= "110000";
        when "0010110101100000" => data <= "110000";
        when "0010110101100001" => data <= "110000";
        when "0010110101100110" => data <= "110000";
        when "0010110101101001" => data <= "110000";
        when "0010110101111101" => data <= "110000";
        when "0010110101111110" => data <= "110000";
        when "0010110101111111" => data <= "110000";
        when "0010110110000000" => data <= "110000";
        when "0010110110001100" => data <= "110000";
        when "0010110110001101" => data <= "001001";
        when "0010110110001110" => data <= "001001";
        when "0010110110001111" => data <= "001001";
        when "0010110110010000" => data <= "001001";
        when "0010110110010001" => data <= "001001";
        when "0010110110010010" => data <= "001001";
        when "0010110110010011" => data <= "001001";
        when "0010110110010100" => data <= "110000";
        when "0010110110011110" => data <= "110000";
        when "0010110110011111" => data <= "110000";
        when "0010111000000000" => data <= "110000";
        when "0010111000000001" => data <= "110000";
        when "0010111000001011" => data <= "110000";
        when "0010111000001100" => data <= "001001";
        when "0010111000001101" => data <= "001001";
        when "0010111000001110" => data <= "001001";
        when "0010111000001111" => data <= "001001";
        when "0010111000010000" => data <= "001001";
        when "0010111000010001" => data <= "001001";
        when "0010111000010010" => data <= "110000";
        when "0010111000011110" => data <= "110000";
        when "0010111000011111" => data <= "110000";
        when "0010111000100100" => data <= "110000";
        when "0010111000100101" => data <= "110000";
        when "0010111000101001" => data <= "110000";
        when "0010111000101010" => data <= "110000";
        when "0010111000101011" => data <= "110000";
        when "0010111000110000" => data <= "110000";
        when "0010111000110001" => data <= "110000";
        when "0010111000110111" => data <= "110000";
        when "0010111000111000" => data <= "110000";
        when "0010111000111001" => data <= "110000";
        when "0010111000111010" => data <= "110000";
        when "0010111000111011" => data <= "110000";
        when "0010111001000000" => data <= "110000";
        when "0010111001000001" => data <= "110000";
        when "0010111001000010" => data <= "110000";
        when "0010111001000011" => data <= "110000";
        when "0010111001000110" => data <= "110000";
        when "0010111001000111" => data <= "110000";
        when "0010111001001010" => data <= "110000";
        when "0010111001001011" => data <= "110000";
        when "0010111001001110" => data <= "110000";
        when "0010111001001111" => data <= "110000";
        when "0010111001010100" => data <= "110000";
        when "0010111001010101" => data <= "110000";
        when "0010111001011001" => data <= "110000";
        when "0010111001011010" => data <= "110000";
        when "0010111001011011" => data <= "110000";
        when "0010111001100000" => data <= "110000";
        when "0010111001100001" => data <= "110000";
        when "0010111001100110" => data <= "110000";
        when "0010111001100111" => data <= "110000";
        when "0010111001101000" => data <= "110000";
        when "0010111001101110" => data <= "110000";
        when "0010111001101111" => data <= "110000";
        when "0010111001110000" => data <= "110000";
        when "0010111001110001" => data <= "110000";
        when "0010111001110101" => data <= "110000";
        when "0010111001110110" => data <= "110000";
        when "0010111001111001" => data <= "110000";
        when "0010111001111010" => data <= "110000";
        when "0010111001111100" => data <= "110000";
        when "0010111001111101" => data <= "110000";
        when "0010111001111111" => data <= "110000";
        when "0010111010000000" => data <= "110000";
        when "0010111010001101" => data <= "110000";
        when "0010111010001110" => data <= "110000";
        when "0010111010001111" => data <= "001001";
        when "0010111010010000" => data <= "001001";
        when "0010111010010001" => data <= "001001";
        when "0010111010010010" => data <= "001001";
        when "0010111010010011" => data <= "001001";
        when "0010111010010100" => data <= "110000";
        when "0010111010011110" => data <= "110000";
        when "0010111010011111" => data <= "110000";
        when "0010111100000000" => data <= "110000";
        when "0010111100000001" => data <= "110000";
        when "0010111100001011" => data <= "110000";
        when "0010111100001100" => data <= "001001";
        when "0010111100001101" => data <= "001001";
        when "0010111100001110" => data <= "001001";
        when "0010111100001111" => data <= "001001";
        when "0010111100010000" => data <= "110000";
        when "0010111100010001" => data <= "110000";
        when "0010111100010100" => data <= "110000";
        when "0010111100011110" => data <= "110000";
        when "0010111100011111" => data <= "110000";
        when "0010111100100100" => data <= "110000";
        when "0010111100100101" => data <= "110000";
        when "0010111100101000" => data <= "110000";
        when "0010111100101100" => data <= "110000";
        when "0010111100110000" => data <= "110000";
        when "0010111100110001" => data <= "110000";
        when "0010111100110011" => data <= "110000";
        when "0010111100110100" => data <= "110000";
        when "0010111100110110" => data <= "110000";
        when "0010111100110111" => data <= "110000";
        when "0010111100111010" => data <= "110000";
        when "0010111100111011" => data <= "110000";
        when "0010111100111111" => data <= "110000";
        when "0010111101000010" => data <= "110000";
        when "0010111101000011" => data <= "110000";
        when "0010111101000110" => data <= "110000";
        when "0010111101000111" => data <= "110000";
        when "0010111101001010" => data <= "110000";
        when "0010111101001011" => data <= "110000";
        when "0010111101001110" => data <= "110000";
        when "0010111101001111" => data <= "110000";
        when "0010111101010100" => data <= "110000";
        when "0010111101010101" => data <= "110000";
        when "0010111101011000" => data <= "110000";
        when "0010111101011100" => data <= "110000";
        when "0010111101100000" => data <= "110000";
        when "0010111101100001" => data <= "110000";
        when "0010111101100110" => data <= "110000";
        when "0010111101100111" => data <= "110000";
        when "0010111101101000" => data <= "110000";
        when "0010111101101001" => data <= "110000";
        when "0010111101101101" => data <= "110000";
        when "0010111101101110" => data <= "110000";
        when "0010111101110010" => data <= "110000";
        when "0010111101110011" => data <= "110000";
        when "0010111101110101" => data <= "110000";
        when "0010111101110110" => data <= "110000";
        when "0010111101111001" => data <= "110000";
        when "0010111101111010" => data <= "110000";
        when "0010111101111100" => data <= "110000";
        when "0010111101111101" => data <= "110000";
        when "0010111110001111" => data <= "110000";
        when "0010111110010000" => data <= "001001";
        when "0010111110010001" => data <= "001001";
        when "0010111110010010" => data <= "001001";
        when "0010111110010011" => data <= "001001";
        when "0010111110010100" => data <= "110000";
        when "0010111110011110" => data <= "110000";
        when "0010111110011111" => data <= "110000";
        when "0011000000000000" => data <= "110000";
        when "0011000000000001" => data <= "110000";
        when "0011000000001011" => data <= "110000";
        when "0011000000001100" => data <= "001001";
        when "0011000000001101" => data <= "001001";
        when "0011000000001110" => data <= "001001";
        when "0011000000001111" => data <= "110000";
        when "0011000000010100" => data <= "110000";
        when "0011000000011110" => data <= "110000";
        when "0011000000011111" => data <= "110000";
        when "0011000000100100" => data <= "110000";
        when "0011000000100101" => data <= "110000";
        when "0011000000100111" => data <= "110000";
        when "0011000000101000" => data <= "110000";
        when "0011000000101100" => data <= "110000";
        when "0011000000101101" => data <= "110000";
        when "0011000000110000" => data <= "110000";
        when "0011000000110001" => data <= "110000";
        when "0011000000110011" => data <= "110000";
        when "0011000000110100" => data <= "110000";
        when "0011000000110110" => data <= "110000";
        when "0011000000110111" => data <= "110000";
        when "0011000000111010" => data <= "110000";
        when "0011000000111011" => data <= "110000";
        when "0011000000111110" => data <= "110000";
        when "0011000000111111" => data <= "110000";
        when "0011000001000010" => data <= "110000";
        when "0011000001000011" => data <= "110000";
        when "0011000001000110" => data <= "110000";
        when "0011000001000111" => data <= "110000";
        when "0011000001001010" => data <= "110000";
        when "0011000001001011" => data <= "110000";
        when "0011000001001110" => data <= "110000";
        when "0011000001001111" => data <= "110000";
        when "0011000001010100" => data <= "110000";
        when "0011000001010101" => data <= "110000";
        when "0011000001010111" => data <= "110000";
        when "0011000001011000" => data <= "110000";
        when "0011000001011100" => data <= "110000";
        when "0011000001011101" => data <= "110000";
        when "0011000001100000" => data <= "110000";
        when "0011000001100001" => data <= "110000";
        when "0011000001100110" => data <= "110000";
        when "0011000001100111" => data <= "110000";
        when "0011000001101010" => data <= "110000";
        when "0011000001101101" => data <= "110000";
        when "0011000001101110" => data <= "110000";
        when "0011000001101111" => data <= "110000";
        when "0011000001110000" => data <= "110000";
        when "0011000001110001" => data <= "110000";
        when "0011000001110010" => data <= "110000";
        when "0011000001110011" => data <= "110000";
        when "0011000001110101" => data <= "110000";
        when "0011000001110110" => data <= "110000";
        when "0011000001111001" => data <= "110000";
        when "0011000001111010" => data <= "110000";
        when "0011000001111101" => data <= "110000";
        when "0011000001111110" => data <= "110000";
        when "0011000001111111" => data <= "110000";
        when "0011000010010000" => data <= "110000";
        when "0011000010010001" => data <= "001001";
        when "0011000010010010" => data <= "001001";
        when "0011000010010011" => data <= "001001";
        when "0011000010010100" => data <= "110000";
        when "0011000010011110" => data <= "110000";
        when "0011000010011111" => data <= "110000";
        when "0011000100000000" => data <= "110000";
        when "0011000100000001" => data <= "110000";
        when "0011000100001011" => data <= "110000";
        when "0011000100001100" => data <= "001001";
        when "0011000100001101" => data <= "001001";
        when "0011000100001110" => data <= "110000";
        when "0011000100010100" => data <= "110000";
        when "0011000100011110" => data <= "110000";
        when "0011000100011111" => data <= "110000";
        when "0011000100100100" => data <= "110000";
        when "0011000100100101" => data <= "110000";
        when "0011000100100111" => data <= "110000";
        when "0011000100101000" => data <= "110000";
        when "0011000100101100" => data <= "110000";
        when "0011000100101101" => data <= "110000";
        when "0011000100110000" => data <= "110000";
        when "0011000100110001" => data <= "110000";
        when "0011000100110011" => data <= "110000";
        when "0011000100110100" => data <= "110000";
        when "0011000100110110" => data <= "110000";
        when "0011000100110111" => data <= "110000";
        when "0011000100111010" => data <= "110000";
        when "0011000100111011" => data <= "110000";
        when "0011000100111110" => data <= "110000";
        when "0011000100111111" => data <= "110000";
        when "0011000101000011" => data <= "110000";
        when "0011000101000100" => data <= "110000";
        when "0011000101000111" => data <= "110000";
        when "0011000101001010" => data <= "110000";
        when "0011000101001110" => data <= "110000";
        when "0011000101001111" => data <= "110000";
        when "0011000101010100" => data <= "110000";
        when "0011000101010101" => data <= "110000";
        when "0011000101010111" => data <= "110000";
        when "0011000101011000" => data <= "110000";
        when "0011000101011100" => data <= "110000";
        when "0011000101011101" => data <= "110000";
        when "0011000101100000" => data <= "110000";
        when "0011000101100001" => data <= "110000";
        when "0011000101100110" => data <= "110000";
        when "0011000101100111" => data <= "110000";
        when "0011000101101010" => data <= "110000";
        when "0011000101101101" => data <= "110000";
        when "0011000101101110" => data <= "110000";
        when "0011000101110110" => data <= "110000";
        when "0011000101111001" => data <= "110000";
        when "0011000101111111" => data <= "110000";
        when "0011000110000000" => data <= "110000";
        when "0011000110001010" => data <= "110000";
        when "0011000110001011" => data <= "110000";
        when "0011000110010001" => data <= "110000";
        when "0011000110010010" => data <= "110000";
        when "0011000110010011" => data <= "001001";
        when "0011000110010100" => data <= "110000";
        when "0011000110011110" => data <= "110000";
        when "0011000110011111" => data <= "110000";
        when "0011001000000000" => data <= "110000";
        when "0011001000000001" => data <= "110000";
        when "0011001000001011" => data <= "110000";
        when "0011001000001100" => data <= "110000";
        when "0011001000001101" => data <= "110000";
        when "0011001000010100" => data <= "110000";
        when "0011001000011110" => data <= "110000";
        when "0011001000011111" => data <= "110000";
        when "0011001000100100" => data <= "110000";
        when "0011001000100101" => data <= "110000";
        when "0011001000101000" => data <= "110000";
        when "0011001000101100" => data <= "110000";
        when "0011001000110000" => data <= "110000";
        when "0011001000110001" => data <= "110000";
        when "0011001000110011" => data <= "110000";
        when "0011001000110100" => data <= "110000";
        when "0011001000110110" => data <= "110000";
        when "0011001000110111" => data <= "110000";
        when "0011001000111010" => data <= "110000";
        when "0011001000111011" => data <= "110000";
        when "0011001000111110" => data <= "110000";
        when "0011001000111111" => data <= "110000";
        when "0011001001000011" => data <= "110000";
        when "0011001001000100" => data <= "110000";
        when "0011001001001000" => data <= "110000";
        when "0011001001001010" => data <= "110000";
        when "0011001001001110" => data <= "110000";
        when "0011001001001111" => data <= "110000";
        when "0011001001010100" => data <= "110000";
        when "0011001001010101" => data <= "110000";
        when "0011001001011000" => data <= "110000";
        when "0011001001011100" => data <= "110000";
        when "0011001001100000" => data <= "110000";
        when "0011001001100001" => data <= "110000";
        when "0011001001100110" => data <= "110000";
        when "0011001001100111" => data <= "110000";
        when "0011001001101010" => data <= "110000";
        when "0011001001101011" => data <= "110000";
        when "0011001001101101" => data <= "110000";
        when "0011001001101110" => data <= "110000";
        when "0011001001110010" => data <= "110000";
        when "0011001001110011" => data <= "110000";
        when "0011001001110111" => data <= "110000";
        when "0011001001111001" => data <= "110000";
        when "0011001001111100" => data <= "110000";
        when "0011001001111101" => data <= "110000";
        when "0011001001111111" => data <= "110000";
        when "0011001010000000" => data <= "110000";
        when "0011001010001010" => data <= "110000";
        when "0011001010001011" => data <= "110000";
        when "0011001010001100" => data <= "110000";
        when "0011001010010011" => data <= "110000";
        when "0011001010010100" => data <= "110000";
        when "0011001010011110" => data <= "110000";
        when "0011001010011111" => data <= "110000";
        when "0011001100000000" => data <= "110000";
        when "0011001100000001" => data <= "110000";
        when "0011001100001011" => data <= "110000";
        when "0011001100010100" => data <= "110000";
        when "0011001100011110" => data <= "110000";
        when "0011001100100100" => data <= "110000";
        when "0011001100101001" => data <= "110000";
        when "0011001100101010" => data <= "110000";
        when "0011001100101011" => data <= "110000";
        when "0011001100101111" => data <= "110000";
        when "0011001100110000" => data <= "110000";
        when "0011001100110001" => data <= "110000";
        when "0011001100110011" => data <= "110000";
        when "0011001100110100" => data <= "110000";
        when "0011001100110111" => data <= "110000";
        when "0011001100111000" => data <= "110000";
        when "0011001100111001" => data <= "110000";
        when "0011001100111010" => data <= "110000";
        when "0011001100111011" => data <= "110000";
        when "0011001100111100" => data <= "110000";
        when "0011001100111111" => data <= "110000";
        when "0011001101000000" => data <= "110000";
        when "0011001101000001" => data <= "110000";
        when "0011001101000010" => data <= "110000";
        when "0011001101000100" => data <= "110000";
        when "0011001101001001" => data <= "110000";
        when "0011001101001010" => data <= "110000";
        when "0011001101001110" => data <= "110000";
        when "0011001101010100" => data <= "110000";
        when "0011001101011001" => data <= "110000";
        when "0011001101011010" => data <= "110000";
        when "0011001101011011" => data <= "110000";
        when "0011001101100000" => data <= "110000";
        when "0011001101100001" => data <= "110000";
        when "0011001101100101" => data <= "110000";
        when "0011001101100110" => data <= "110000";
        when "0011001101100111" => data <= "110000";
        when "0011001101101010" => data <= "110000";
        when "0011001101101011" => data <= "110000";
        when "0011001101101110" => data <= "110000";
        when "0011001101101111" => data <= "110000";
        when "0011001101110000" => data <= "110000";
        when "0011001101110001" => data <= "110000";
        when "0011001101110010" => data <= "110000";
        when "0011001101111000" => data <= "110000";
        when "0011001101111001" => data <= "110000";
        when "0011001101111100" => data <= "110000";
        when "0011001101111101" => data <= "110000";
        when "0011001101111110" => data <= "110000";
        when "0011001101111111" => data <= "110000";
        when "0011001110001010" => data <= "110000";
        when "0011001110001100" => data <= "110000";
        when "0011001110001101" => data <= "110000";
        when "0011001110010100" => data <= "110000";
        when "0011001110011110" => data <= "110000";
        when "0011001110011111" => data <= "110000";
        when "0011010000000000" => data <= "110000";
        when "0011010000000001" => data <= "110000";
        when "0011010000001001" => data <= "110000";
        when "0011010000001010" => data <= "110000";
        when "0011010000001011" => data <= "110000";
        when "0011010000010100" => data <= "110000";
        when "0011010001000110" => data <= "110000";
        when "0011010001000111" => data <= "110000";
        when "0011010001001001" => data <= "110000";
        when "0011010001001010" => data <= "110000";
        when "0011010001110101" => data <= "110000";
        when "0011010001110110" => data <= "110000";
        when "0011010001111000" => data <= "110000";
        when "0011010001111001" => data <= "110000";
        when "0011010010001010" => data <= "110000";
        when "0011010010001101" => data <= "110000";
        when "0011010010001110" => data <= "110000";
        when "0011010010010100" => data <= "110000";
        when "0011010010010101" => data <= "110000";
        when "0011010010010110" => data <= "110000";
        when "0011010010011110" => data <= "110000";
        when "0011010010011111" => data <= "110000";
        when "0011010100000000" => data <= "110000";
        when "0011010100000001" => data <= "110000";
        when "0011010100001000" => data <= "110000";
        when "0011010100001001" => data <= "001001";
        when "0011010100001010" => data <= "001001";
        when "0011010100001011" => data <= "110000";
        when "0011010100010100" => data <= "110000";
        when "0011010101000110" => data <= "110000";
        when "0011010101000111" => data <= "110000";
        when "0011010101001000" => data <= "110000";
        when "0011010101001001" => data <= "110000";
        when "0011010101110101" => data <= "110000";
        when "0011010101110110" => data <= "110000";
        when "0011010101110111" => data <= "110000";
        when "0011010101111000" => data <= "110000";
        when "0011010110001010" => data <= "110000";
        when "0011010110001110" => data <= "110000";
        when "0011010110010100" => data <= "110000";
        when "0011010110010101" => data <= "001001";
        when "0011010110010110" => data <= "001001";
        when "0011010110010111" => data <= "110000";
        when "0011010110011110" => data <= "110000";
        when "0011010110011111" => data <= "110000";
        when "0011011000000000" => data <= "110000";
        when "0011011000000001" => data <= "110000";
        when "0011011000000111" => data <= "110000";
        when "0011011000001000" => data <= "001001";
        when "0011011000001001" => data <= "001001";
        when "0011011000001010" => data <= "001001";
        when "0011011000001011" => data <= "110000";
        when "0011011000010001" => data <= "110000";
        when "0011011000010010" => data <= "110000";
        when "0011011000010011" => data <= "110000";
        when "0011011000010100" => data <= "110000";
        when "0011011010001010" => data <= "110000";
        when "0011011010001110" => data <= "110000";
        when "0011011010001111" => data <= "110000";
        when "0011011010010100" => data <= "110000";
        when "0011011010010101" => data <= "001001";
        when "0011011010010110" => data <= "001001";
        when "0011011010010111" => data <= "001001";
        when "0011011010011000" => data <= "110000";
        when "0011011010011110" => data <= "110000";
        when "0011011010011111" => data <= "110000";
        when "0011011100000000" => data <= "110000";
        when "0011011100000001" => data <= "110000";
        when "0011011100000101" => data <= "110000";
        when "0011011100000110" => data <= "110000";
        when "0011011100000111" => data <= "001001";
        when "0011011100001000" => data <= "001001";
        when "0011011100001001" => data <= "001001";
        when "0011011100001010" => data <= "001001";
        when "0011011100001011" => data <= "110000";
        when "0011011100010000" => data <= "110000";
        when "0011011100010001" => data <= "110000";
        when "0011011100010010" => data <= "110000";
        when "0011011100010011" => data <= "110000";
        when "0011011100010100" => data <= "110000";
        when "0011011110001010" => data <= "110000";
        when "0011011110001111" => data <= "110000";
        when "0011011110010100" => data <= "110000";
        when "0011011110010101" => data <= "001001";
        when "0011011110010110" => data <= "001001";
        when "0011011110010111" => data <= "001001";
        when "0011011110011000" => data <= "001001";
        when "0011011110011001" => data <= "110000";
        when "0011011110011010" => data <= "110000";
        when "0011011110011110" => data <= "110000";
        when "0011011110011111" => data <= "110000";
        when "0011100000000000" => data <= "110000";
        when "0011100000000001" => data <= "110000";
        when "0011100000000100" => data <= "110000";
        when "0011100000000101" => data <= "001001";
        when "0011100000000110" => data <= "001001";
        when "0011100000000111" => data <= "001001";
        when "0011100000001000" => data <= "001001";
        when "0011100000001001" => data <= "001001";
        when "0011100000001010" => data <= "001001";
        when "0011100000001011" => data <= "110000";
        when "0011100000001111" => data <= "110000";
        when "0011100000010000" => data <= "110000";
        when "0011100000010001" => data <= "110000";
        when "0011100000010010" => data <= "110000";
        when "0011100000010011" => data <= "110000";
        when "0011100000010100" => data <= "110000";
        when "0011100000110100" => data <= "111111";
        when "0011100000110101" => data <= "111111";
        when "0011100000110110" => data <= "111111";
        when "0011100000110111" => data <= "111111";
        when "0011100001010011" => data <= "111111";
        when "0011100001010100" => data <= "111111";
        when "0011100001010101" => data <= "111111";
        when "0011100001010110" => data <= "111111";
        when "0011100001011001" => data <= "111111";
        when "0011100001101001" => data <= "111111";
        when "0011100010001010" => data <= "110000";
        when "0011100010010100" => data <= "110000";
        when "0011100010010101" => data <= "001001";
        when "0011100010010110" => data <= "001001";
        when "0011100010010111" => data <= "001001";
        when "0011100010011000" => data <= "001001";
        when "0011100010011001" => data <= "001001";
        when "0011100010011010" => data <= "001001";
        when "0011100010011011" => data <= "110000";
        when "0011100010011110" => data <= "110000";
        when "0011100010011111" => data <= "110000";
        when "0011100100000000" => data <= "110000";
        when "0011100100000001" => data <= "110000";
        when "0011100100000011" => data <= "110000";
        when "0011100100000100" => data <= "001001";
        when "0011100100000101" => data <= "001001";
        when "0011100100000110" => data <= "001001";
        when "0011100100000111" => data <= "001001";
        when "0011100100001000" => data <= "001001";
        when "0011100100001001" => data <= "001001";
        when "0011100100001010" => data <= "001001";
        when "0011100100001011" => data <= "110000";
        when "0011100100001111" => data <= "110000";
        when "0011100100010000" => data <= "110000";
        when "0011100100010001" => data <= "110000";
        when "0011100100010010" => data <= "110000";
        when "0011100100010011" => data <= "110000";
        when "0011100100010100" => data <= "110000";
        when "0011100100110100" => data <= "111111";
        when "0011100100111000" => data <= "111111";
        when "0011100101010010" => data <= "111111";
        when "0011100101011001" => data <= "111111";
        when "0011100101101001" => data <= "111111";
        when "0011100110001010" => data <= "110000";
        when "0011100110010100" => data <= "110000";
        when "0011100110010101" => data <= "001001";
        when "0011100110010110" => data <= "001001";
        when "0011100110010111" => data <= "001001";
        when "0011100110011000" => data <= "001001";
        when "0011100110011001" => data <= "001001";
        when "0011100110011010" => data <= "001001";
        when "0011100110011011" => data <= "001001";
        when "0011100110011100" => data <= "110000";
        when "0011100110011110" => data <= "110000";
        when "0011100110011111" => data <= "110000";
        when "0011101000000000" => data <= "110000";
        when "0011101000000001" => data <= "110000";
        when "0011101000000010" => data <= "110000";
        when "0011101000000011" => data <= "001001";
        when "0011101000000100" => data <= "001001";
        when "0011101000000101" => data <= "001001";
        when "0011101000000110" => data <= "001001";
        when "0011101000000111" => data <= "001001";
        when "0011101000001000" => data <= "001001";
        when "0011101000001001" => data <= "001001";
        when "0011101000001010" => data <= "001001";
        when "0011101000001011" => data <= "110000";
        when "0011101000001111" => data <= "110000";
        when "0011101000010000" => data <= "110000";
        when "0011101000010001" => data <= "110000";
        when "0011101000010010" => data <= "110000";
        when "0011101000010011" => data <= "110000";
        when "0011101000010100" => data <= "110000";
        when "0011101000110100" => data <= "111111";
        when "0011101000111000" => data <= "111111";
        when "0011101000111010" => data <= "111111";
        when "0011101000111100" => data <= "111111";
        when "0011101000111101" => data <= "111111";
        when "0011101001000000" => data <= "111111";
        when "0011101001000001" => data <= "111111";
        when "0011101001000010" => data <= "111111";
        when "0011101001000110" => data <= "111111";
        when "0011101001000111" => data <= "111111";
        when "0011101001001000" => data <= "111111";
        when "0011101001001001" => data <= "111111";
        when "0011101001001100" => data <= "111111";
        when "0011101001001101" => data <= "111111";
        when "0011101001001110" => data <= "111111";
        when "0011101001001111" => data <= "111111";
        when "0011101001010010" => data <= "111111";
        when "0011101001011000" => data <= "111111";
        when "0011101001011001" => data <= "111111";
        when "0011101001011010" => data <= "111111";
        when "0011101001011011" => data <= "111111";
        when "0011101001011110" => data <= "111111";
        when "0011101001011111" => data <= "111111";
        when "0011101001100000" => data <= "111111";
        when "0011101001100011" => data <= "111111";
        when "0011101001100101" => data <= "111111";
        when "0011101001100110" => data <= "111111";
        when "0011101001101000" => data <= "111111";
        when "0011101001101001" => data <= "111111";
        when "0011101001101010" => data <= "111111";
        when "0011101001101011" => data <= "111111";
        when "0011101010001010" => data <= "110000";
        when "0011101010010100" => data <= "110000";
        when "0011101010010101" => data <= "001001";
        when "0011101010010110" => data <= "001001";
        when "0011101010010111" => data <= "001001";
        when "0011101010011000" => data <= "001001";
        when "0011101010011001" => data <= "001001";
        when "0011101010011010" => data <= "001001";
        when "0011101010011011" => data <= "001001";
        when "0011101010011100" => data <= "001001";
        when "0011101010011101" => data <= "110000";
        when "0011101010011110" => data <= "110000";
        when "0011101010011111" => data <= "110000";
        when "0011101100000000" => data <= "110000";
        when "0011101100000001" => data <= "110000";
        when "0011101100000010" => data <= "001001";
        when "0011101100000011" => data <= "001001";
        when "0011101100000100" => data <= "001001";
        when "0011101100000101" => data <= "001001";
        when "0011101100000110" => data <= "001001";
        when "0011101100000111" => data <= "001001";
        when "0011101100001000" => data <= "001001";
        when "0011101100001001" => data <= "001001";
        when "0011101100001010" => data <= "001001";
        when "0011101100001011" => data <= "110000";
        when "0011101100001111" => data <= "110000";
        when "0011101100010000" => data <= "110000";
        when "0011101100010001" => data <= "110000";
        when "0011101100010010" => data <= "110000";
        when "0011101100010011" => data <= "110000";
        when "0011101100010100" => data <= "110000";
        when "0011101100110100" => data <= "111111";
        when "0011101100111000" => data <= "111111";
        when "0011101100111010" => data <= "111111";
        when "0011101100111011" => data <= "111111";
        when "0011101100111111" => data <= "111111";
        when "0011101101000011" => data <= "111111";
        when "0011101101000101" => data <= "111111";
        when "0011101101001011" => data <= "111111";
        when "0011101101010011" => data <= "111111";
        when "0011101101010100" => data <= "111111";
        when "0011101101010101" => data <= "111111";
        when "0011101101011001" => data <= "111111";
        when "0011101101100001" => data <= "111111";
        when "0011101101100011" => data <= "111111";
        when "0011101101100100" => data <= "111111";
        when "0011101101101001" => data <= "111111";
        when "0011101110000111" => data <= "110000";
        when "0011101110001000" => data <= "110000";
        when "0011101110001010" => data <= "110000";
        when "0011101110010100" => data <= "110000";
        when "0011101110010101" => data <= "001001";
        when "0011101110010110" => data <= "001001";
        when "0011101110010111" => data <= "001001";
        when "0011101110011000" => data <= "001001";
        when "0011101110011001" => data <= "001001";
        when "0011101110011010" => data <= "001001";
        when "0011101110011011" => data <= "001001";
        when "0011101110011100" => data <= "001001";
        when "0011101110011101" => data <= "001001";
        when "0011101110011110" => data <= "110000";
        when "0011101110011111" => data <= "110000";
        when "0011110000000000" => data <= "110000";
        when "0011110000000001" => data <= "110000";
        when "0011110000000010" => data <= "110000";
        when "0011110000000011" => data <= "001001";
        when "0011110000000100" => data <= "001001";
        when "0011110000000101" => data <= "001001";
        when "0011110000000110" => data <= "001001";
        when "0011110000000111" => data <= "001001";
        when "0011110000001000" => data <= "001001";
        when "0011110000001001" => data <= "001001";
        when "0011110000001010" => data <= "001001";
        when "0011110000001011" => data <= "110000";
        when "0011110000001111" => data <= "110000";
        when "0011110000010000" => data <= "110000";
        when "0011110000010001" => data <= "110000";
        when "0011110000010010" => data <= "110000";
        when "0011110000010011" => data <= "110000";
        when "0011110000010100" => data <= "110000";
        when "0011110000110100" => data <= "111111";
        when "0011110000110101" => data <= "111111";
        when "0011110000110110" => data <= "111111";
        when "0011110000110111" => data <= "111111";
        when "0011110000111010" => data <= "111111";
        when "0011110000111111" => data <= "111111";
        when "0011110001000000" => data <= "111111";
        when "0011110001000001" => data <= "111111";
        when "0011110001000010" => data <= "111111";
        when "0011110001000011" => data <= "111111";
        when "0011110001000110" => data <= "111111";
        when "0011110001000111" => data <= "111111";
        when "0011110001001000" => data <= "111111";
        when "0011110001001100" => data <= "111111";
        when "0011110001001101" => data <= "111111";
        when "0011110001001110" => data <= "111111";
        when "0011110001010110" => data <= "111111";
        when "0011110001011001" => data <= "111111";
        when "0011110001011110" => data <= "111111";
        when "0011110001011111" => data <= "111111";
        when "0011110001100000" => data <= "111111";
        when "0011110001100001" => data <= "111111";
        when "0011110001100011" => data <= "111111";
        when "0011110001101001" => data <= "111111";
        when "0011110010000110" => data <= "110000";
        when "0011110010000111" => data <= "110000";
        when "0011110010001000" => data <= "110000";
        when "0011110010001001" => data <= "110000";
        when "0011110010001010" => data <= "110000";
        when "0011110010010100" => data <= "110000";
        when "0011110010010101" => data <= "001001";
        when "0011110010010110" => data <= "001001";
        when "0011110010010111" => data <= "001001";
        when "0011110010011000" => data <= "001001";
        when "0011110010011001" => data <= "001001";
        when "0011110010011010" => data <= "001001";
        when "0011110010011011" => data <= "001001";
        when "0011110010011100" => data <= "001001";
        when "0011110010011101" => data <= "110000";
        when "0011110010011110" => data <= "110000";
        when "0011110010011111" => data <= "110000";
        when "0011110100000000" => data <= "110000";
        when "0011110100000001" => data <= "110000";
        when "0011110100000011" => data <= "110000";
        when "0011110100000100" => data <= "001001";
        when "0011110100000101" => data <= "001001";
        when "0011110100000110" => data <= "001001";
        when "0011110100000111" => data <= "001001";
        when "0011110100001000" => data <= "001001";
        when "0011110100001001" => data <= "001001";
        when "0011110100001010" => data <= "001001";
        when "0011110100001011" => data <= "110000";
        when "0011110100001111" => data <= "110000";
        when "0011110100010000" => data <= "110000";
        when "0011110100010001" => data <= "110000";
        when "0011110100010010" => data <= "110000";
        when "0011110100010011" => data <= "110000";
        when "0011110100010100" => data <= "110000";
        when "0011110100110100" => data <= "111111";
        when "0011110100111010" => data <= "111111";
        when "0011110100111111" => data <= "111111";
        when "0011110101001001" => data <= "111111";
        when "0011110101001111" => data <= "111111";
        when "0011110101010110" => data <= "111111";
        when "0011110101011001" => data <= "111111";
        when "0011110101011101" => data <= "111111";
        when "0011110101100001" => data <= "111111";
        when "0011110101100011" => data <= "111111";
        when "0011110101101001" => data <= "111111";
        when "0011110110000101" => data <= "110000";
        when "0011110110000110" => data <= "110000";
        when "0011110110001010" => data <= "110000";
        when "0011110110010100" => data <= "110000";
        when "0011110110010101" => data <= "001001";
        when "0011110110010110" => data <= "001001";
        when "0011110110010111" => data <= "001001";
        when "0011110110011000" => data <= "001001";
        when "0011110110011001" => data <= "001001";
        when "0011110110011010" => data <= "001001";
        when "0011110110011011" => data <= "001001";
        when "0011110110011100" => data <= "110000";
        when "0011110110011110" => data <= "110000";
        when "0011110110011111" => data <= "110000";
        when "0011111000000000" => data <= "110000";
        when "0011111000000001" => data <= "110000";
        when "0011111000000100" => data <= "110000";
        when "0011111000000101" => data <= "001001";
        when "0011111000000110" => data <= "001001";
        when "0011111000000111" => data <= "001001";
        when "0011111000001000" => data <= "001001";
        when "0011111000001001" => data <= "001001";
        when "0011111000001010" => data <= "001001";
        when "0011111000001011" => data <= "110000";
        when "0011111000010000" => data <= "110000";
        when "0011111000010001" => data <= "110000";
        when "0011111000010010" => data <= "110000";
        when "0011111000010011" => data <= "110000";
        when "0011111000010100" => data <= "110000";
        when "0011111000110100" => data <= "111111";
        when "0011111000111010" => data <= "111111";
        when "0011111001000000" => data <= "111111";
        when "0011111001000001" => data <= "111111";
        when "0011111001000010" => data <= "111111";
        when "0011111001000101" => data <= "111111";
        when "0011111001000110" => data <= "111111";
        when "0011111001000111" => data <= "111111";
        when "0011111001001000" => data <= "111111";
        when "0011111001001011" => data <= "111111";
        when "0011111001001100" => data <= "111111";
        when "0011111001001101" => data <= "111111";
        when "0011111001001110" => data <= "111111";
        when "0011111001010010" => data <= "111111";
        when "0011111001010011" => data <= "111111";
        when "0011111001010100" => data <= "111111";
        when "0011111001010101" => data <= "111111";
        when "0011111001011010" => data <= "111111";
        when "0011111001011011" => data <= "111111";
        when "0011111001011110" => data <= "111111";
        when "0011111001011111" => data <= "111111";
        when "0011111001100000" => data <= "111111";
        when "0011111001100001" => data <= "111111";
        when "0011111001100011" => data <= "111111";
        when "0011111001101010" => data <= "111111";
        when "0011111001101011" => data <= "111111";
        when "0011111010000101" => data <= "110000";
        when "0011111010001010" => data <= "110000";
        when "0011111010010100" => data <= "110000";
        when "0011111010010101" => data <= "001001";
        when "0011111010010110" => data <= "001001";
        when "0011111010010111" => data <= "001001";
        when "0011111010011000" => data <= "001001";
        when "0011111010011001" => data <= "001001";
        when "0011111010011010" => data <= "001001";
        when "0011111010011011" => data <= "110000";
        when "0011111010011110" => data <= "110000";
        when "0011111010011111" => data <= "110000";
        when "0011111100000000" => data <= "110000";
        when "0011111100000001" => data <= "110000";
        when "0011111100000101" => data <= "110000";
        when "0011111100000110" => data <= "110000";
        when "0011111100000111" => data <= "001001";
        when "0011111100001000" => data <= "001001";
        when "0011111100001001" => data <= "001001";
        when "0011111100001010" => data <= "001001";
        when "0011111100001011" => data <= "110000";
        when "0011111100010000" => data <= "110000";
        when "0011111100010001" => data <= "110000";
        when "0011111100010010" => data <= "110000";
        when "0011111100010011" => data <= "110000";
        when "0011111100010100" => data <= "110000";
        when "0011111110000101" => data <= "110000";
        when "0011111110001010" => data <= "110000";
        when "0011111110010100" => data <= "110000";
        when "0011111110010101" => data <= "001001";
        when "0011111110010110" => data <= "001001";
        when "0011111110010111" => data <= "001001";
        when "0011111110011000" => data <= "001001";
        when "0011111110011001" => data <= "110000";
        when "0011111110011010" => data <= "110000";
        when "0011111110011110" => data <= "110000";
        when "0011111110011111" => data <= "110000";
        when "0100000000000000" => data <= "110000";
        when "0100000000000001" => data <= "110000";
        when "0100000000000111" => data <= "110000";
        when "0100000000001000" => data <= "001001";
        when "0100000000001001" => data <= "001001";
        when "0100000000001010" => data <= "001001";
        when "0100000000001011" => data <= "110000";
        when "0100000000010100" => data <= "110000";
        when "0100000010000101" => data <= "110000";
        when "0100000010001010" => data <= "110000";
        when "0100000010010100" => data <= "110000";
        when "0100000010010101" => data <= "001001";
        when "0100000010010110" => data <= "001001";
        when "0100000010010111" => data <= "001001";
        when "0100000010011000" => data <= "110000";
        when "0100000010011110" => data <= "110000";
        when "0100000010011111" => data <= "110000";
        when "0100000100000000" => data <= "110000";
        when "0100000100000001" => data <= "110000";
        when "0100000100001000" => data <= "110000";
        when "0100000100001001" => data <= "001001";
        when "0100000100001010" => data <= "001001";
        when "0100000100001011" => data <= "110000";
        when "0100000110000101" => data <= "110000";
        when "0100000110000110" => data <= "110000";
        when "0100000110001010" => data <= "110000";
        when "0100000110010100" => data <= "110000";
        when "0100000110010101" => data <= "001001";
        when "0100000110010110" => data <= "001001";
        when "0100000110010111" => data <= "110000";
        when "0100000110011110" => data <= "110000";
        when "0100000110011111" => data <= "110000";
        when "0100001000000000" => data <= "110000";
        when "0100001000000001" => data <= "110000";
        when "0100001000001001" => data <= "110000";
        when "0100001000001010" => data <= "110000";
        when "0100001000001011" => data <= "110000";
        when "0100001010000110" => data <= "110000";
        when "0100001010000111" => data <= "110000";
        when "0100001010001000" => data <= "110000";
        when "0100001010001001" => data <= "110000";
        when "0100001010001010" => data <= "110000";
        when "0100001010010100" => data <= "110000";
        when "0100001010010101" => data <= "001001";
        when "0100001010010110" => data <= "110000";
        when "0100001010011110" => data <= "110000";
        when "0100001010011111" => data <= "110000";
        when "0100001100000000" => data <= "110000";
        when "0100001100000001" => data <= "110000";
        when "0100001100001011" => data <= "110000";
        when "0100001110010100" => data <= "110000";
        when "0100001110010101" => data <= "110000";
        when "0100001110011110" => data <= "110000";
        when "0100001110011111" => data <= "110000";
        when "0100010000000000" => data <= "110000";
        when "0100010000000001" => data <= "110000";
        when "0100010000001011" => data <= "110000";
        when "0100010000001100" => data <= "110000";
        when "0100010010010011" => data <= "110000";
        when "0100010010010100" => data <= "110000";
        when "0100010010011110" => data <= "110000";
        when "0100010010011111" => data <= "110000";
        when "0100010100000000" => data <= "110000";
        when "0100010100000001" => data <= "110000";
        when "0100010100001011" => data <= "110000";
        when "0100010100001100" => data <= "001001";
        when "0100010100001101" => data <= "110000";
        when "0100010100001110" => data <= "110000";
        when "0100010110010010" => data <= "110000";
        when "0100010110010011" => data <= "001001";
        when "0100010110010100" => data <= "110000";
        when "0100010110011110" => data <= "110000";
        when "0100010110011111" => data <= "110000";
        when "0100011000000000" => data <= "110000";
        when "0100011000000001" => data <= "110000";
        when "0100011000001011" => data <= "110000";
        when "0100011000001100" => data <= "001001";
        when "0100011000001101" => data <= "001001";
        when "0100011000001110" => data <= "001001";
        when "0100011000001111" => data <= "110000";
        when "0100011010010000" => data <= "110000";
        when "0100011010010001" => data <= "110000";
        when "0100011010010010" => data <= "001001";
        when "0100011010010011" => data <= "001001";
        when "0100011010010100" => data <= "110000";
        when "0100011010011110" => data <= "110000";
        when "0100011010011111" => data <= "110000";
        when "0100011100000000" => data <= "110000";
        when "0100011100000001" => data <= "110000";
        when "0100011100001011" => data <= "110000";
        when "0100011100001100" => data <= "001001";
        when "0100011100001101" => data <= "001001";
        when "0100011100001110" => data <= "001001";
        when "0100011100001111" => data <= "001001";
        when "0100011100010000" => data <= "110000";
        when "0100011110001111" => data <= "110000";
        when "0100011110010000" => data <= "001001";
        when "0100011110010001" => data <= "001001";
        when "0100011110010010" => data <= "001001";
        when "0100011110010011" => data <= "001001";
        when "0100011110010100" => data <= "110000";
        when "0100011110011110" => data <= "110000";
        when "0100011110011111" => data <= "110000";
        when "0100100000000000" => data <= "110000";
        when "0100100000000001" => data <= "110000";
        when "0100100000001011" => data <= "110000";
        when "0100100000001100" => data <= "001001";
        when "0100100000001101" => data <= "001001";
        when "0100100000001110" => data <= "001001";
        when "0100100000001111" => data <= "001001";
        when "0100100000010000" => data <= "001001";
        when "0100100000010001" => data <= "110000";
        when "0100100000010010" => data <= "110000";
        when "0100100010001110" => data <= "110000";
        when "0100100010001111" => data <= "001001";
        when "0100100010010000" => data <= "001001";
        when "0100100010010001" => data <= "001001";
        when "0100100010010010" => data <= "001001";
        when "0100100010010011" => data <= "001001";
        when "0100100010010100" => data <= "110000";
        when "0100100010011110" => data <= "110000";
        when "0100100010011111" => data <= "110000";
        when "0100100100000000" => data <= "110000";
        when "0100100100000001" => data <= "110000";
        when "0100100100001011" => data <= "110000";
        when "0100100100001100" => data <= "001001";
        when "0100100100001101" => data <= "001001";
        when "0100100100001110" => data <= "001001";
        when "0100100100001111" => data <= "001001";
        when "0100100100010000" => data <= "001001";
        when "0100100100010001" => data <= "001001";
        when "0100100100010010" => data <= "001001";
        when "0100100100010011" => data <= "110000";
        when "0100100110001100" => data <= "110000";
        when "0100100110001101" => data <= "110000";
        when "0100100110001110" => data <= "001001";
        when "0100100110001111" => data <= "001001";
        when "0100100110010000" => data <= "001001";
        when "0100100110010001" => data <= "001001";
        when "0100100110010010" => data <= "001001";
        when "0100100110010011" => data <= "001001";
        when "0100100110010100" => data <= "110000";
        when "0100100110011110" => data <= "110000";
        when "0100100110011111" => data <= "110000";
        when "0100101000000000" => data <= "110000";
        when "0100101000000001" => data <= "110000";
        when "0100101000001011" => data <= "110000";
        when "0100101000001100" => data <= "001001";
        when "0100101000001101" => data <= "001001";
        when "0100101000001110" => data <= "001001";
        when "0100101000001111" => data <= "001001";
        when "0100101000010000" => data <= "001001";
        when "0100101000010001" => data <= "001001";
        when "0100101000010010" => data <= "001001";
        when "0100101000010011" => data <= "001001";
        when "0100101000010100" => data <= "110000";
        when "0100101010001011" => data <= "110000";
        when "0100101010001100" => data <= "001001";
        when "0100101010001101" => data <= "001001";
        when "0100101010001110" => data <= "001001";
        when "0100101010001111" => data <= "001001";
        when "0100101010010000" => data <= "001001";
        when "0100101010010001" => data <= "001001";
        when "0100101010010010" => data <= "001001";
        when "0100101010010011" => data <= "001001";
        when "0100101010010100" => data <= "110000";
        when "0100101010011110" => data <= "110000";
        when "0100101010011111" => data <= "110000";
        when "0100101100000000" => data <= "110000";
        when "0100101100000001" => data <= "110000";
        when "0100101100001011" => data <= "110000";
        when "0100101100001100" => data <= "001001";
        when "0100101100001101" => data <= "001001";
        when "0100101100001110" => data <= "001001";
        when "0100101100001111" => data <= "001001";
        when "0100101100010000" => data <= "001001";
        when "0100101100010001" => data <= "001001";
        when "0100101100010010" => data <= "001001";
        when "0100101100010011" => data <= "001001";
        when "0100101100010100" => data <= "001001";
        when "0100101100010101" => data <= "110000";
        when "0100101100010110" => data <= "110000";
        when "0100101110001010" => data <= "110000";
        when "0100101110001011" => data <= "001001";
        when "0100101110001100" => data <= "001001";
        when "0100101110001101" => data <= "001001";
        when "0100101110001110" => data <= "001001";
        when "0100101110001111" => data <= "001001";
        when "0100101110010000" => data <= "001001";
        when "0100101110010001" => data <= "001001";
        when "0100101110010010" => data <= "001001";
        when "0100101110010011" => data <= "001001";
        when "0100101110010100" => data <= "110000";
        when "0100101110011110" => data <= "110000";
        when "0100101110011111" => data <= "110000";
        when "0100110000000000" => data <= "110000";
        when "0100110000000001" => data <= "110000";
        when "0100110000001011" => data <= "110000";
        when "0100110000001100" => data <= "001001";
        when "0100110000001101" => data <= "001001";
        when "0100110000001110" => data <= "001001";
        when "0100110000001111" => data <= "001001";
        when "0100110000010000" => data <= "001001";
        when "0100110000010001" => data <= "001001";
        when "0100110000010010" => data <= "001001";
        when "0100110000010011" => data <= "001001";
        when "0100110000010100" => data <= "001001";
        when "0100110000010101" => data <= "001001";
        when "0100110000010110" => data <= "001001";
        when "0100110000010111" => data <= "110000";
        when "0100110010001000" => data <= "110000";
        when "0100110010001001" => data <= "110000";
        when "0100110010001010" => data <= "001001";
        when "0100110010001011" => data <= "001001";
        when "0100110010001100" => data <= "001001";
        when "0100110010001101" => data <= "001001";
        when "0100110010001110" => data <= "001001";
        when "0100110010001111" => data <= "001001";
        when "0100110010010000" => data <= "001001";
        when "0100110010010001" => data <= "001001";
        when "0100110010010010" => data <= "001001";
        when "0100110010010011" => data <= "001001";
        when "0100110010010100" => data <= "110000";
        when "0100110010011110" => data <= "110000";
        when "0100110010011111" => data <= "110000";
        when "0100110100000000" => data <= "110000";
        when "0100110100000001" => data <= "110000";
        when "0100110100001011" => data <= "110000";
        when "0100110100001100" => data <= "001001";
        when "0100110100001101" => data <= "001001";
        when "0100110100001110" => data <= "001001";
        when "0100110100001111" => data <= "001001";
        when "0100110100010000" => data <= "001001";
        when "0100110100010001" => data <= "001001";
        when "0100110100010010" => data <= "001001";
        when "0100110100010011" => data <= "001001";
        when "0100110100010100" => data <= "001001";
        when "0100110100010101" => data <= "001001";
        when "0100110100010110" => data <= "001001";
        when "0100110100010111" => data <= "001001";
        when "0100110100011000" => data <= "110000";
        when "0100110110000111" => data <= "110000";
        when "0100110110001000" => data <= "001001";
        when "0100110110001001" => data <= "001001";
        when "0100110110001010" => data <= "001001";
        when "0100110110001011" => data <= "001001";
        when "0100110110001100" => data <= "001001";
        when "0100110110001101" => data <= "001001";
        when "0100110110001110" => data <= "001001";
        when "0100110110001111" => data <= "001001";
        when "0100110110010000" => data <= "001001";
        when "0100110110010001" => data <= "001001";
        when "0100110110010010" => data <= "001001";
        when "0100110110010011" => data <= "001001";
        when "0100110110010100" => data <= "110000";
        when "0100110110011110" => data <= "110000";
        when "0100110110011111" => data <= "110000";
        when "0100111000000000" => data <= "110000";
        when "0100111000000001" => data <= "110000";
        when "0100111000001011" => data <= "110000";
        when "0100111000001100" => data <= "001001";
        when "0100111000001101" => data <= "001001";
        when "0100111000001110" => data <= "001001";
        when "0100111000001111" => data <= "001001";
        when "0100111000010000" => data <= "001001";
        when "0100111000010001" => data <= "001001";
        when "0100111000010010" => data <= "001001";
        when "0100111000010011" => data <= "001001";
        when "0100111000010100" => data <= "001001";
        when "0100111000010101" => data <= "001001";
        when "0100111000010110" => data <= "001001";
        when "0100111000010111" => data <= "001001";
        when "0100111000011000" => data <= "001001";
        when "0100111000011001" => data <= "110000";
        when "0100111000011010" => data <= "110000";
        when "0100111010000110" => data <= "110000";
        when "0100111010000111" => data <= "001001";
        when "0100111010001000" => data <= "001001";
        when "0100111010001001" => data <= "001001";
        when "0100111010001010" => data <= "001001";
        when "0100111010001011" => data <= "001001";
        when "0100111010001100" => data <= "001001";
        when "0100111010001101" => data <= "001001";
        when "0100111010001110" => data <= "001001";
        when "0100111010001111" => data <= "001001";
        when "0100111010010000" => data <= "001001";
        when "0100111010010001" => data <= "001001";
        when "0100111010010010" => data <= "001001";
        when "0100111010010011" => data <= "001001";
        when "0100111010010100" => data <= "110000";
        when "0100111010011110" => data <= "110000";
        when "0100111010011111" => data <= "110000";
        when "0100111100000000" => data <= "110000";
        when "0100111100000001" => data <= "110000";
        when "0100111100001011" => data <= "110000";
        when "0100111100001100" => data <= "001001";
        when "0100111100001101" => data <= "001001";
        when "0100111100001110" => data <= "001001";
        when "0100111100001111" => data <= "001001";
        when "0100111100010000" => data <= "001001";
        when "0100111100010001" => data <= "001001";
        when "0100111100010010" => data <= "001001";
        when "0100111100010011" => data <= "001001";
        when "0100111100010100" => data <= "001001";
        when "0100111100010101" => data <= "001001";
        when "0100111100010110" => data <= "001001";
        when "0100111100010111" => data <= "001001";
        when "0100111100011000" => data <= "001001";
        when "0100111100011001" => data <= "001001";
        when "0100111100011010" => data <= "001001";
        when "0100111100011011" => data <= "110000";
        when "0100111110000100" => data <= "110000";
        when "0100111110000101" => data <= "110000";
        when "0100111110000110" => data <= "001001";
        when "0100111110000111" => data <= "001001";
        when "0100111110001000" => data <= "001001";
        when "0100111110001001" => data <= "001001";
        when "0100111110001010" => data <= "001001";
        when "0100111110001011" => data <= "001001";
        when "0100111110001100" => data <= "001001";
        when "0100111110001101" => data <= "001001";
        when "0100111110001110" => data <= "001001";
        when "0100111110001111" => data <= "001001";
        when "0100111110010000" => data <= "001001";
        when "0100111110010001" => data <= "001001";
        when "0100111110010010" => data <= "001001";
        when "0100111110010011" => data <= "001001";
        when "0100111110010100" => data <= "110000";
        when "0100111110011110" => data <= "110000";
        when "0100111110011111" => data <= "110000";
        when "0101000000000000" => data <= "110000";
        when "0101000000000001" => data <= "110000";
        when "0101000000001011" => data <= "110000";
        when "0101000000001100" => data <= "001001";
        when "0101000000001101" => data <= "001001";
        when "0101000000001110" => data <= "001001";
        when "0101000000001111" => data <= "001001";
        when "0101000000010000" => data <= "001001";
        when "0101000000010001" => data <= "001001";
        when "0101000000010010" => data <= "001001";
        when "0101000000010011" => data <= "001001";
        when "0101000000010100" => data <= "001001";
        when "0101000000010101" => data <= "001001";
        when "0101000000010110" => data <= "001001";
        when "0101000000010111" => data <= "001001";
        when "0101000000011000" => data <= "001001";
        when "0101000000011001" => data <= "001001";
        when "0101000000011010" => data <= "001001";
        when "0101000000011011" => data <= "001001";
        when "0101000000011100" => data <= "110000";
        when "0101000010000011" => data <= "110000";
        when "0101000010000100" => data <= "001001";
        when "0101000010000101" => data <= "001001";
        when "0101000010000110" => data <= "001001";
        when "0101000010000111" => data <= "001001";
        when "0101000010001000" => data <= "001001";
        when "0101000010001001" => data <= "001001";
        when "0101000010001010" => data <= "001001";
        when "0101000010001011" => data <= "001001";
        when "0101000010001100" => data <= "001001";
        when "0101000010001101" => data <= "001001";
        when "0101000010001110" => data <= "001001";
        when "0101000010001111" => data <= "001001";
        when "0101000010010000" => data <= "001001";
        when "0101000010010001" => data <= "001001";
        when "0101000010010010" => data <= "001001";
        when "0101000010010011" => data <= "001001";
        when "0101000010010100" => data <= "110000";
        when "0101000010011110" => data <= "110000";
        when "0101000010011111" => data <= "110000";
        when "0101000100000000" => data <= "110000";
        when "0101000100000001" => data <= "110000";
        when "0101000100001011" => data <= "110000";
        when "0101000100001100" => data <= "001001";
        when "0101000100001101" => data <= "001001";
        when "0101000100001110" => data <= "001001";
        when "0101000100001111" => data <= "001001";
        when "0101000100010000" => data <= "001001";
        when "0101000100010001" => data <= "001001";
        when "0101000100010010" => data <= "001001";
        when "0101000100010011" => data <= "001001";
        when "0101000100010100" => data <= "001001";
        when "0101000100010101" => data <= "001001";
        when "0101000100010110" => data <= "001001";
        when "0101000100010111" => data <= "001001";
        when "0101000100011000" => data <= "001001";
        when "0101000100011001" => data <= "001001";
        when "0101000100011010" => data <= "001001";
        when "0101000100011011" => data <= "001001";
        when "0101000100011100" => data <= "001001";
        when "0101000100011101" => data <= "110000";
        when "0101000100011110" => data <= "110000";
        when "0101000110000010" => data <= "110000";
        when "0101000110000011" => data <= "001001";
        when "0101000110000100" => data <= "001001";
        when "0101000110000101" => data <= "001001";
        when "0101000110000110" => data <= "001001";
        when "0101000110000111" => data <= "001001";
        when "0101000110001000" => data <= "001001";
        when "0101000110001001" => data <= "001001";
        when "0101000110001010" => data <= "001001";
        when "0101000110001011" => data <= "001001";
        when "0101000110001100" => data <= "001001";
        when "0101000110001101" => data <= "001001";
        when "0101000110001110" => data <= "001001";
        when "0101000110001111" => data <= "001001";
        when "0101000110010000" => data <= "001001";
        when "0101000110010001" => data <= "001001";
        when "0101000110010010" => data <= "001001";
        when "0101000110010011" => data <= "001001";
        when "0101000110010100" => data <= "110000";
        when "0101000110011110" => data <= "110000";
        when "0101000110011111" => data <= "110000";
        when "0101001000000000" => data <= "110000";
        when "0101001000000001" => data <= "110000";
        when "0101001000001011" => data <= "110000";
        when "0101001000001100" => data <= "001001";
        when "0101001000001101" => data <= "001001";
        when "0101001000001110" => data <= "001001";
        when "0101001000001111" => data <= "001001";
        when "0101001000010000" => data <= "001001";
        when "0101001000010001" => data <= "001001";
        when "0101001000010010" => data <= "001001";
        when "0101001000010011" => data <= "001001";
        when "0101001000010100" => data <= "001001";
        when "0101001000010101" => data <= "001001";
        when "0101001000010110" => data <= "001001";
        when "0101001000010111" => data <= "001001";
        when "0101001000011000" => data <= "001001";
        when "0101001000011001" => data <= "001001";
        when "0101001000011010" => data <= "001001";
        when "0101001000011011" => data <= "001001";
        when "0101001000011100" => data <= "001001";
        when "0101001000011101" => data <= "001001";
        when "0101001000011110" => data <= "001001";
        when "0101001000011111" => data <= "110000";
        when "0101001010000001" => data <= "110000";
        when "0101001010000010" => data <= "001001";
        when "0101001010000011" => data <= "001001";
        when "0101001010000100" => data <= "001001";
        when "0101001010000101" => data <= "001001";
        when "0101001010000110" => data <= "001001";
        when "0101001010000111" => data <= "001001";
        when "0101001010001000" => data <= "001001";
        when "0101001010001001" => data <= "001001";
        when "0101001010001010" => data <= "001001";
        when "0101001010001011" => data <= "001001";
        when "0101001010001100" => data <= "001001";
        when "0101001010001101" => data <= "001001";
        when "0101001010001110" => data <= "001001";
        when "0101001010001111" => data <= "001001";
        when "0101001010010000" => data <= "001001";
        when "0101001010010001" => data <= "001001";
        when "0101001010010010" => data <= "001001";
        when "0101001010010011" => data <= "001001";
        when "0101001010010100" => data <= "110000";
        when "0101001010011110" => data <= "110000";
        when "0101001010011111" => data <= "110000";
        when "0101001100000000" => data <= "110000";
        when "0101001100000001" => data <= "110000";
        when "0101001100001011" => data <= "110000";
        when "0101001100001100" => data <= "001001";
        when "0101001100001101" => data <= "001001";
        when "0101001100001110" => data <= "001001";
        when "0101001100001111" => data <= "001001";
        when "0101001100010000" => data <= "001001";
        when "0101001100010001" => data <= "001001";
        when "0101001100010010" => data <= "001001";
        when "0101001100010011" => data <= "001001";
        when "0101001100010100" => data <= "001001";
        when "0101001100010101" => data <= "001001";
        when "0101001100010110" => data <= "001001";
        when "0101001100010111" => data <= "001001";
        when "0101001100011000" => data <= "001001";
        when "0101001100011001" => data <= "001001";
        when "0101001100011010" => data <= "001001";
        when "0101001100011011" => data <= "001001";
        when "0101001100011100" => data <= "001001";
        when "0101001100011101" => data <= "001001";
        when "0101001100011110" => data <= "001001";
        when "0101001100011111" => data <= "001001";
        when "0101001100100000" => data <= "110000";
        when "0101001101111111" => data <= "110000";
        when "0101001110000000" => data <= "110000";
        when "0101001110000001" => data <= "001001";
        when "0101001110000010" => data <= "001001";
        when "0101001110000011" => data <= "001001";
        when "0101001110000100" => data <= "001001";
        when "0101001110000101" => data <= "001001";
        when "0101001110000110" => data <= "001001";
        when "0101001110000111" => data <= "001001";
        when "0101001110001000" => data <= "001001";
        when "0101001110001001" => data <= "001001";
        when "0101001110001010" => data <= "001001";
        when "0101001110001011" => data <= "001001";
        when "0101001110001100" => data <= "001001";
        when "0101001110001101" => data <= "001001";
        when "0101001110001110" => data <= "001001";
        when "0101001110001111" => data <= "001001";
        when "0101001110010000" => data <= "001001";
        when "0101001110010001" => data <= "001001";
        when "0101001110010010" => data <= "001001";
        when "0101001110010011" => data <= "001001";
        when "0101001110010100" => data <= "110000";
        when "0101001110011110" => data <= "110000";
        when "0101001110011111" => data <= "110000";
        when "0101010000000000" => data <= "110000";
        when "0101010000000001" => data <= "110000";
        when "0101010000001011" => data <= "110000";
        when "0101010000001100" => data <= "001001";
        when "0101010000001101" => data <= "001001";
        when "0101010000001110" => data <= "001001";
        when "0101010000001111" => data <= "001001";
        when "0101010000010000" => data <= "001001";
        when "0101010000010001" => data <= "001001";
        when "0101010000010010" => data <= "001001";
        when "0101010000010011" => data <= "001001";
        when "0101010000010100" => data <= "001001";
        when "0101010000010101" => data <= "001001";
        when "0101010000010110" => data <= "001001";
        when "0101010000010111" => data <= "001001";
        when "0101010000011000" => data <= "001001";
        when "0101010000011001" => data <= "001001";
        when "0101010000011010" => data <= "001001";
        when "0101010000011011" => data <= "001001";
        when "0101010000011100" => data <= "001001";
        when "0101010000011101" => data <= "001001";
        when "0101010000011110" => data <= "001001";
        when "0101010000011111" => data <= "001001";
        when "0101010000100000" => data <= "001001";
        when "0101010000100001" => data <= "110000";
        when "0101010000100010" => data <= "110000";
        when "0101010001111110" => data <= "110000";
        when "0101010001111111" => data <= "001001";
        when "0101010010000000" => data <= "001001";
        when "0101010010000001" => data <= "001001";
        when "0101010010000010" => data <= "001001";
        when "0101010010000011" => data <= "001001";
        when "0101010010000100" => data <= "001001";
        when "0101010010000101" => data <= "001001";
        when "0101010010000110" => data <= "001001";
        when "0101010010000111" => data <= "001001";
        when "0101010010001000" => data <= "001001";
        when "0101010010001001" => data <= "001001";
        when "0101010010001010" => data <= "001001";
        when "0101010010001011" => data <= "001001";
        when "0101010010001100" => data <= "001001";
        when "0101010010001101" => data <= "001001";
        when "0101010010001110" => data <= "001001";
        when "0101010010001111" => data <= "001001";
        when "0101010010010000" => data <= "001001";
        when "0101010010010001" => data <= "001001";
        when "0101010010010010" => data <= "001001";
        when "0101010010010011" => data <= "001001";
        when "0101010010010100" => data <= "110000";
        when "0101010010011110" => data <= "110000";
        when "0101010010011111" => data <= "110000";
        when "0101010100000000" => data <= "110000";
        when "0101010100000001" => data <= "110000";
        when "0101010100001011" => data <= "110000";
        when "0101010100001100" => data <= "001001";
        when "0101010100001101" => data <= "001001";
        when "0101010100001110" => data <= "001001";
        when "0101010100001111" => data <= "001001";
        when "0101010100010000" => data <= "001001";
        when "0101010100010001" => data <= "001001";
        when "0101010100010010" => data <= "001001";
        when "0101010100010011" => data <= "001001";
        when "0101010100010100" => data <= "001001";
        when "0101010100010101" => data <= "001001";
        when "0101010100010110" => data <= "001001";
        when "0101010100010111" => data <= "001001";
        when "0101010100011000" => data <= "001001";
        when "0101010100011001" => data <= "001001";
        when "0101010100011010" => data <= "001001";
        when "0101010100011011" => data <= "001001";
        when "0101010100011100" => data <= "001001";
        when "0101010100011101" => data <= "001001";
        when "0101010100011110" => data <= "001001";
        when "0101010100011111" => data <= "001001";
        when "0101010100100000" => data <= "001001";
        when "0101010100100001" => data <= "001001";
        when "0101010100100010" => data <= "001001";
        when "0101010100100011" => data <= "110000";
        when "0101010101111101" => data <= "110000";
        when "0101010101111110" => data <= "001001";
        when "0101010101111111" => data <= "001001";
        when "0101010110000000" => data <= "001001";
        when "0101010110000001" => data <= "001001";
        when "0101010110000010" => data <= "001001";
        when "0101010110000011" => data <= "001001";
        when "0101010110000100" => data <= "001001";
        when "0101010110000101" => data <= "001001";
        when "0101010110000110" => data <= "001001";
        when "0101010110000111" => data <= "001001";
        when "0101010110001000" => data <= "001001";
        when "0101010110001001" => data <= "001001";
        when "0101010110001010" => data <= "001001";
        when "0101010110001011" => data <= "001001";
        when "0101010110001100" => data <= "001001";
        when "0101010110001101" => data <= "001001";
        when "0101010110001110" => data <= "001001";
        when "0101010110001111" => data <= "001001";
        when "0101010110010000" => data <= "001001";
        when "0101010110010001" => data <= "001001";
        when "0101010110010010" => data <= "001001";
        when "0101010110010011" => data <= "001001";
        when "0101010110010100" => data <= "110000";
        when "0101010110011110" => data <= "110000";
        when "0101010110011111" => data <= "110000";
        when "0101011000000000" => data <= "110000";
        when "0101011000000001" => data <= "110000";
        when "0101011000001011" => data <= "110000";
        when "0101011000001100" => data <= "001001";
        when "0101011000001101" => data <= "001001";
        when "0101011000001110" => data <= "001001";
        when "0101011000001111" => data <= "001001";
        when "0101011000010000" => data <= "001001";
        when "0101011000010001" => data <= "001001";
        when "0101011000010010" => data <= "001001";
        when "0101011000010011" => data <= "001001";
        when "0101011000010100" => data <= "001001";
        when "0101011000010101" => data <= "001001";
        when "0101011000010110" => data <= "001001";
        when "0101011000010111" => data <= "001001";
        when "0101011000011000" => data <= "001001";
        when "0101011000011001" => data <= "001001";
        when "0101011000011010" => data <= "001001";
        when "0101011000011011" => data <= "001001";
        when "0101011000011100" => data <= "001001";
        when "0101011000011101" => data <= "001001";
        when "0101011000011110" => data <= "001001";
        when "0101011000011111" => data <= "001001";
        when "0101011000100000" => data <= "001001";
        when "0101011000100001" => data <= "001001";
        when "0101011000100010" => data <= "001001";
        when "0101011000100011" => data <= "001001";
        when "0101011000100100" => data <= "110000";
        when "0101011001111011" => data <= "110000";
        when "0101011001111100" => data <= "110000";
        when "0101011001111101" => data <= "001001";
        when "0101011001111110" => data <= "001001";
        when "0101011001111111" => data <= "001001";
        when "0101011010000000" => data <= "001001";
        when "0101011010000001" => data <= "001001";
        when "0101011010000010" => data <= "001001";
        when "0101011010000011" => data <= "001001";
        when "0101011010000100" => data <= "001001";
        when "0101011010000101" => data <= "001001";
        when "0101011010000110" => data <= "001001";
        when "0101011010000111" => data <= "001001";
        when "0101011010001000" => data <= "001001";
        when "0101011010001001" => data <= "001001";
        when "0101011010001010" => data <= "001001";
        when "0101011010001011" => data <= "001001";
        when "0101011010001100" => data <= "001001";
        when "0101011010001101" => data <= "001001";
        when "0101011010001110" => data <= "001001";
        when "0101011010001111" => data <= "001001";
        when "0101011010010000" => data <= "001001";
        when "0101011010010001" => data <= "001001";
        when "0101011010010010" => data <= "001001";
        when "0101011010010011" => data <= "001001";
        when "0101011010010100" => data <= "110000";
        when "0101011010011110" => data <= "110000";
        when "0101011010011111" => data <= "110000";
        when "0101011100000000" => data <= "110000";
        when "0101011100000001" => data <= "110000";
        when "0101011100001011" => data <= "110000";
        when "0101011100001100" => data <= "001001";
        when "0101011100001101" => data <= "001001";
        when "0101011100001110" => data <= "001001";
        when "0101011100001111" => data <= "001001";
        when "0101011100010000" => data <= "001001";
        when "0101011100010001" => data <= "001001";
        when "0101011100010010" => data <= "001001";
        when "0101011100010011" => data <= "001001";
        when "0101011100010100" => data <= "001001";
        when "0101011100010101" => data <= "001001";
        when "0101011100010110" => data <= "001001";
        when "0101011100010111" => data <= "001001";
        when "0101011100011000" => data <= "001001";
        when "0101011100011001" => data <= "001001";
        when "0101011100011010" => data <= "001001";
        when "0101011100011011" => data <= "001001";
        when "0101011100011100" => data <= "001001";
        when "0101011100011101" => data <= "001001";
        when "0101011100011110" => data <= "001001";
        when "0101011100011111" => data <= "001001";
        when "0101011100100000" => data <= "001001";
        when "0101011100100001" => data <= "001001";
        when "0101011100100010" => data <= "001001";
        when "0101011100100011" => data <= "001001";
        when "0101011100100100" => data <= "001001";
        when "0101011100100101" => data <= "110000";
        when "0101011100100110" => data <= "110000";
        when "0101011101111010" => data <= "110000";
        when "0101011101111011" => data <= "001001";
        when "0101011101111100" => data <= "001001";
        when "0101011101111101" => data <= "001001";
        when "0101011101111110" => data <= "001001";
        when "0101011101111111" => data <= "001001";
        when "0101011110000000" => data <= "001001";
        when "0101011110000001" => data <= "001001";
        when "0101011110000010" => data <= "001001";
        when "0101011110000011" => data <= "001001";
        when "0101011110000100" => data <= "001001";
        when "0101011110000101" => data <= "001001";
        when "0101011110000110" => data <= "001001";
        when "0101011110000111" => data <= "001001";
        when "0101011110001000" => data <= "001001";
        when "0101011110001001" => data <= "001001";
        when "0101011110001010" => data <= "001001";
        when "0101011110001011" => data <= "001001";
        when "0101011110001100" => data <= "001001";
        when "0101011110001101" => data <= "001001";
        when "0101011110001110" => data <= "001001";
        when "0101011110001111" => data <= "001001";
        when "0101011110010000" => data <= "001001";
        when "0101011110010001" => data <= "001001";
        when "0101011110010010" => data <= "001001";
        when "0101011110010011" => data <= "001001";
        when "0101011110010100" => data <= "110000";
        when "0101011110011110" => data <= "110000";
        when "0101011110011111" => data <= "110000";
        when "0101100000000000" => data <= "110000";
        when "0101100000000001" => data <= "110000";
        when "0101100000001011" => data <= "110000";
        when "0101100000001100" => data <= "001001";
        when "0101100000001101" => data <= "001001";
        when "0101100000001110" => data <= "001001";
        when "0101100000001111" => data <= "001001";
        when "0101100000010000" => data <= "001001";
        when "0101100000010001" => data <= "001001";
        when "0101100000010010" => data <= "001001";
        when "0101100000010011" => data <= "001001";
        when "0101100000010100" => data <= "001001";
        when "0101100000010101" => data <= "001001";
        when "0101100000010110" => data <= "001001";
        when "0101100000010111" => data <= "001001";
        when "0101100000011000" => data <= "001001";
        when "0101100000011001" => data <= "001001";
        when "0101100000011010" => data <= "001001";
        when "0101100000011011" => data <= "001001";
        when "0101100000011100" => data <= "001001";
        when "0101100000011101" => data <= "001001";
        when "0101100000011110" => data <= "001001";
        when "0101100000011111" => data <= "001001";
        when "0101100000100000" => data <= "001001";
        when "0101100000100001" => data <= "001001";
        when "0101100000100010" => data <= "001001";
        when "0101100000100011" => data <= "001001";
        when "0101100000100100" => data <= "001001";
        when "0101100000100101" => data <= "001001";
        when "0101100000100110" => data <= "001001";
        when "0101100000100111" => data <= "110000";
        when "0101100001111001" => data <= "110000";
        when "0101100001111010" => data <= "001001";
        when "0101100001111011" => data <= "001001";
        when "0101100001111100" => data <= "001001";
        when "0101100001111101" => data <= "001001";
        when "0101100001111110" => data <= "001001";
        when "0101100001111111" => data <= "001001";
        when "0101100010000000" => data <= "001001";
        when "0101100010000001" => data <= "001001";
        when "0101100010000010" => data <= "001001";
        when "0101100010000011" => data <= "001001";
        when "0101100010000100" => data <= "001001";
        when "0101100010000101" => data <= "001001";
        when "0101100010000110" => data <= "001001";
        when "0101100010000111" => data <= "001001";
        when "0101100010001000" => data <= "001001";
        when "0101100010001001" => data <= "001001";
        when "0101100010001010" => data <= "001001";
        when "0101100010001011" => data <= "001001";
        when "0101100010001100" => data <= "001001";
        when "0101100010001101" => data <= "001001";
        when "0101100010001110" => data <= "001001";
        when "0101100010001111" => data <= "001001";
        when "0101100010010000" => data <= "001001";
        when "0101100010010001" => data <= "001001";
        when "0101100010010010" => data <= "001001";
        when "0101100010010011" => data <= "001001";
        when "0101100010010100" => data <= "110000";
        when "0101100010011110" => data <= "110000";
        when "0101100010011111" => data <= "110000";
        when "0101100100000000" => data <= "110000";
        when "0101100100000001" => data <= "110000";
        when "0101100100001011" => data <= "110000";
        when "0101100100001100" => data <= "110000";
        when "0101100100001101" => data <= "001001";
        when "0101100100001110" => data <= "001001";
        when "0101100100001111" => data <= "001001";
        when "0101100100010000" => data <= "001001";
        when "0101100100010001" => data <= "001001";
        when "0101100100010010" => data <= "001001";
        when "0101100100010011" => data <= "001001";
        when "0101100100010100" => data <= "001001";
        when "0101100100010101" => data <= "001001";
        when "0101100100010110" => data <= "001001";
        when "0101100100010111" => data <= "001001";
        when "0101100100011000" => data <= "001001";
        when "0101100100011001" => data <= "001001";
        when "0101100100011010" => data <= "001001";
        when "0101100100011011" => data <= "001001";
        when "0101100100011100" => data <= "001001";
        when "0101100100011101" => data <= "001001";
        when "0101100100011110" => data <= "001001";
        when "0101100100011111" => data <= "001001";
        when "0101100100100000" => data <= "001001";
        when "0101100100100001" => data <= "001001";
        when "0101100100100010" => data <= "001001";
        when "0101100100100011" => data <= "001001";
        when "0101100100100100" => data <= "001001";
        when "0101100100100101" => data <= "001001";
        when "0101100100100110" => data <= "001001";
        when "0101100100100111" => data <= "001001";
        when "0101100100101000" => data <= "110000";
        when "0101100101110111" => data <= "110000";
        when "0101100101111000" => data <= "110000";
        when "0101100101111001" => data <= "001001";
        when "0101100101111010" => data <= "001001";
        when "0101100101111011" => data <= "001001";
        when "0101100101111100" => data <= "001001";
        when "0101100101111101" => data <= "001001";
        when "0101100101111110" => data <= "001001";
        when "0101100101111111" => data <= "001001";
        when "0101100110000000" => data <= "001001";
        when "0101100110000001" => data <= "001001";
        when "0101100110000010" => data <= "001001";
        when "0101100110000011" => data <= "001001";
        when "0101100110000100" => data <= "001001";
        when "0101100110000101" => data <= "001001";
        when "0101100110000110" => data <= "001001";
        when "0101100110000111" => data <= "001001";
        when "0101100110001000" => data <= "001001";
        when "0101100110001001" => data <= "001001";
        when "0101100110001010" => data <= "001001";
        when "0101100110001011" => data <= "001001";
        when "0101100110001100" => data <= "001001";
        when "0101100110001101" => data <= "001001";
        when "0101100110001110" => data <= "001001";
        when "0101100110001111" => data <= "001001";
        when "0101100110010000" => data <= "001001";
        when "0101100110010001" => data <= "001001";
        when "0101100110010010" => data <= "001001";
        when "0101100110010011" => data <= "110000";
        when "0101100110010100" => data <= "110000";
        when "0101100110011110" => data <= "110000";
        when "0101100110011111" => data <= "110000";
        when "0101101000000000" => data <= "110000";
        when "0101101000000001" => data <= "110000";
        when "0101101000001101" => data <= "110000";
        when "0101101000001110" => data <= "110000";
        when "0101101000001111" => data <= "110000";
        when "0101101000010000" => data <= "001001";
        when "0101101000010001" => data <= "001001";
        when "0101101000010010" => data <= "001001";
        when "0101101000010011" => data <= "001001";
        when "0101101000010100" => data <= "001001";
        when "0101101000010101" => data <= "001001";
        when "0101101000010110" => data <= "001001";
        when "0101101000010111" => data <= "001001";
        when "0101101000011000" => data <= "001001";
        when "0101101000011001" => data <= "001001";
        when "0101101000011010" => data <= "001001";
        when "0101101000011011" => data <= "001001";
        when "0101101000011100" => data <= "001001";
        when "0101101000011101" => data <= "001001";
        when "0101101000011110" => data <= "001001";
        when "0101101000011111" => data <= "001001";
        when "0101101000100000" => data <= "001001";
        when "0101101000100001" => data <= "001001";
        when "0101101000100010" => data <= "001001";
        when "0101101000100011" => data <= "001001";
        when "0101101000100100" => data <= "001001";
        when "0101101000100101" => data <= "001001";
        when "0101101000100110" => data <= "001001";
        when "0101101000100111" => data <= "001001";
        when "0101101000101000" => data <= "001001";
        when "0101101000101001" => data <= "110000";
        when "0101101001001010" => data <= "110000";
        when "0101101001001011" => data <= "110000";
        when "0101101001001100" => data <= "110000";
        when "0101101001001101" => data <= "110000";
        when "0101101001001110" => data <= "110000";
        when "0101101001001111" => data <= "110000";
        when "0101101001010000" => data <= "110000";
        when "0101101001010001" => data <= "110000";
        when "0101101001010010" => data <= "110000";
        when "0101101001010011" => data <= "110000";
        when "0101101001010100" => data <= "110000";
        when "0101101001010101" => data <= "110000";
        when "0101101001010110" => data <= "110000";
        when "0101101001010111" => data <= "110000";
        when "0101101001011000" => data <= "110000";
        when "0101101001110110" => data <= "110000";
        when "0101101001110111" => data <= "001001";
        when "0101101001111000" => data <= "001001";
        when "0101101001111001" => data <= "001001";
        when "0101101001111010" => data <= "001001";
        when "0101101001111011" => data <= "001001";
        when "0101101001111100" => data <= "001001";
        when "0101101001111101" => data <= "001001";
        when "0101101001111110" => data <= "001001";
        when "0101101001111111" => data <= "001001";
        when "0101101010000000" => data <= "001001";
        when "0101101010000001" => data <= "001001";
        when "0101101010000010" => data <= "001001";
        when "0101101010000011" => data <= "001001";
        when "0101101010000100" => data <= "001001";
        when "0101101010000101" => data <= "001001";
        when "0101101010000110" => data <= "001001";
        when "0101101010000111" => data <= "001001";
        when "0101101010001000" => data <= "001001";
        when "0101101010001001" => data <= "001001";
        when "0101101010001010" => data <= "001001";
        when "0101101010001011" => data <= "001001";
        when "0101101010001100" => data <= "001001";
        when "0101101010001101" => data <= "001001";
        when "0101101010001110" => data <= "001001";
        when "0101101010001111" => data <= "001001";
        when "0101101010010000" => data <= "001001";
        when "0101101010010001" => data <= "110000";
        when "0101101010010010" => data <= "110000";
        when "0101101010011110" => data <= "110000";
        when "0101101010011111" => data <= "110000";
        when "0101101100000000" => data <= "110000";
        when "0101101100000001" => data <= "110000";
        when "0101101100010000" => data <= "110000";
        when "0101101100010001" => data <= "110000";
        when "0101101100010010" => data <= "001001";
        when "0101101100010011" => data <= "001001";
        when "0101101100010100" => data <= "001001";
        when "0101101100010101" => data <= "001001";
        when "0101101100010110" => data <= "001001";
        when "0101101100010111" => data <= "001001";
        when "0101101100011000" => data <= "001001";
        when "0101101100011001" => data <= "001001";
        when "0101101100011010" => data <= "001001";
        when "0101101100011011" => data <= "001001";
        when "0101101100011100" => data <= "001001";
        when "0101101100011101" => data <= "001001";
        when "0101101100011110" => data <= "001001";
        when "0101101100011111" => data <= "001001";
        when "0101101100100000" => data <= "001001";
        when "0101101100100001" => data <= "001001";
        when "0101101100100010" => data <= "001001";
        when "0101101100100011" => data <= "001001";
        when "0101101100100100" => data <= "001001";
        when "0101101100100101" => data <= "001001";
        when "0101101100100110" => data <= "001001";
        when "0101101100100111" => data <= "001001";
        when "0101101100101000" => data <= "001001";
        when "0101101100101001" => data <= "001001";
        when "0101101100101010" => data <= "110000";
        when "0101101100101011" => data <= "110000";
        when "0101101101001010" => data <= "110000";
        when "0101101101011000" => data <= "110000";
        when "0101101101110101" => data <= "110000";
        when "0101101101110110" => data <= "001001";
        when "0101101101110111" => data <= "001001";
        when "0101101101111000" => data <= "001001";
        when "0101101101111001" => data <= "001001";
        when "0101101101111010" => data <= "001001";
        when "0101101101111011" => data <= "001001";
        when "0101101101111100" => data <= "001001";
        when "0101101101111101" => data <= "001001";
        when "0101101101111110" => data <= "001001";
        when "0101101101111111" => data <= "001001";
        when "0101101110000000" => data <= "001001";
        when "0101101110000001" => data <= "001001";
        when "0101101110000010" => data <= "001001";
        when "0101101110000011" => data <= "001001";
        when "0101101110000100" => data <= "001001";
        when "0101101110000101" => data <= "001001";
        when "0101101110000110" => data <= "001001";
        when "0101101110000111" => data <= "001001";
        when "0101101110001000" => data <= "001001";
        when "0101101110001001" => data <= "001001";
        when "0101101110001010" => data <= "001001";
        when "0101101110001011" => data <= "001001";
        when "0101101110001100" => data <= "001001";
        when "0101101110001101" => data <= "001001";
        when "0101101110001110" => data <= "110000";
        when "0101101110001111" => data <= "110000";
        when "0101101110010000" => data <= "110000";
        when "0101101110011110" => data <= "110000";
        when "0101101110011111" => data <= "110000";
        when "0101110000000000" => data <= "110000";
        when "0101110000000001" => data <= "110000";
        when "0101110000010010" => data <= "110000";
        when "0101110000010011" => data <= "110000";
        when "0101110000010100" => data <= "001001";
        when "0101110000010101" => data <= "001001";
        when "0101110000010110" => data <= "001001";
        when "0101110000010111" => data <= "001001";
        when "0101110000011000" => data <= "001001";
        when "0101110000011001" => data <= "001001";
        when "0101110000011010" => data <= "001001";
        when "0101110000011011" => data <= "001001";
        when "0101110000011100" => data <= "001001";
        when "0101110000011101" => data <= "001001";
        when "0101110000011110" => data <= "001001";
        when "0101110000011111" => data <= "001001";
        when "0101110000100000" => data <= "001001";
        when "0101110000100001" => data <= "001001";
        when "0101110000100010" => data <= "001001";
        when "0101110000100011" => data <= "001001";
        when "0101110000100100" => data <= "001001";
        when "0101110000100101" => data <= "001001";
        when "0101110000100110" => data <= "001001";
        when "0101110000100111" => data <= "001001";
        when "0101110000101000" => data <= "001001";
        when "0101110000101001" => data <= "001001";
        when "0101110000101010" => data <= "001001";
        when "0101110000101011" => data <= "001001";
        when "0101110000101100" => data <= "110000";
        when "0101110001001010" => data <= "110000";
        when "0101110001001011" => data <= "110000";
        when "0101110001001100" => data <= "110000";
        when "0101110001001101" => data <= "110000";
        when "0101110001001110" => data <= "110000";
        when "0101110001001111" => data <= "110000";
        when "0101110001010000" => data <= "110000";
        when "0101110001010001" => data <= "110000";
        when "0101110001010010" => data <= "110000";
        when "0101110001010011" => data <= "110000";
        when "0101110001010100" => data <= "110000";
        when "0101110001010101" => data <= "110000";
        when "0101110001010110" => data <= "110000";
        when "0101110001010111" => data <= "110000";
        when "0101110001011000" => data <= "110000";
        when "0101110001110011" => data <= "110000";
        when "0101110001110100" => data <= "110000";
        when "0101110001110101" => data <= "001001";
        when "0101110001110110" => data <= "001001";
        when "0101110001110111" => data <= "001001";
        when "0101110001111000" => data <= "001001";
        when "0101110001111001" => data <= "001001";
        when "0101110001111010" => data <= "001001";
        when "0101110001111011" => data <= "001001";
        when "0101110001111100" => data <= "001001";
        when "0101110001111101" => data <= "001001";
        when "0101110001111110" => data <= "001001";
        when "0101110001111111" => data <= "001001";
        when "0101110010000000" => data <= "001001";
        when "0101110010000001" => data <= "001001";
        when "0101110010000010" => data <= "001001";
        when "0101110010000011" => data <= "001001";
        when "0101110010000100" => data <= "001001";
        when "0101110010000101" => data <= "001001";
        when "0101110010000110" => data <= "001001";
        when "0101110010000111" => data <= "001001";
        when "0101110010001000" => data <= "001001";
        when "0101110010001001" => data <= "001001";
        when "0101110010001010" => data <= "001001";
        when "0101110010001011" => data <= "001001";
        when "0101110010001100" => data <= "110000";
        when "0101110010001101" => data <= "110000";
        when "0101110010011110" => data <= "110000";
        when "0101110010011111" => data <= "110000";
        when "0101110100000000" => data <= "110000";
        when "0101110100000001" => data <= "110000";
        when "0101110100010100" => data <= "110000";
        when "0101110100010101" => data <= "110000";
        when "0101110100010110" => data <= "001001";
        when "0101110100010111" => data <= "001001";
        when "0101110100011000" => data <= "001001";
        when "0101110100011001" => data <= "001001";
        when "0101110100011010" => data <= "001001";
        when "0101110100011011" => data <= "001001";
        when "0101110100011100" => data <= "001001";
        when "0101110100011101" => data <= "001001";
        when "0101110100011110" => data <= "001001";
        when "0101110100011111" => data <= "001001";
        when "0101110100100000" => data <= "001001";
        when "0101110100100001" => data <= "001001";
        when "0101110100100010" => data <= "001001";
        when "0101110100100011" => data <= "001001";
        when "0101110100100100" => data <= "001001";
        when "0101110100100101" => data <= "001001";
        when "0101110100100110" => data <= "001001";
        when "0101110100100111" => data <= "001001";
        when "0101110100101000" => data <= "001001";
        when "0101110100101001" => data <= "001001";
        when "0101110100101010" => data <= "001001";
        when "0101110100101011" => data <= "001001";
        when "0101110100101100" => data <= "001001";
        when "0101110100101101" => data <= "110000";
        when "0101110101001010" => data <= "110000";
        when "0101110101011000" => data <= "110000";
        when "0101110101110010" => data <= "110000";
        when "0101110101110011" => data <= "001001";
        when "0101110101110100" => data <= "001001";
        when "0101110101110101" => data <= "001001";
        when "0101110101110110" => data <= "001001";
        when "0101110101110111" => data <= "001001";
        when "0101110101111000" => data <= "001001";
        when "0101110101111001" => data <= "001001";
        when "0101110101111010" => data <= "001001";
        when "0101110101111011" => data <= "001001";
        when "0101110101111100" => data <= "001001";
        when "0101110101111101" => data <= "001001";
        when "0101110101111110" => data <= "001001";
        when "0101110101111111" => data <= "001001";
        when "0101110110000000" => data <= "001001";
        when "0101110110000001" => data <= "001001";
        when "0101110110000010" => data <= "001001";
        when "0101110110000011" => data <= "001001";
        when "0101110110000100" => data <= "001001";
        when "0101110110000101" => data <= "001001";
        when "0101110110000110" => data <= "001001";
        when "0101110110000111" => data <= "001001";
        when "0101110110001000" => data <= "001001";
        when "0101110110001001" => data <= "001001";
        when "0101110110001010" => data <= "110000";
        when "0101110110001011" => data <= "110000";
        when "0101110110011110" => data <= "110000";
        when "0101110110011111" => data <= "110000";
        when "0101111000000000" => data <= "110000";
        when "0101111000000001" => data <= "110000";
        when "0101111000010110" => data <= "110000";
        when "0101111000010111" => data <= "110000";
        when "0101111000011000" => data <= "110000";
        when "0101111000011001" => data <= "001001";
        when "0101111000011010" => data <= "001001";
        when "0101111000011011" => data <= "001001";
        when "0101111000011100" => data <= "001001";
        when "0101111000011101" => data <= "001001";
        when "0101111000011110" => data <= "001001";
        when "0101111000011111" => data <= "001001";
        when "0101111000100000" => data <= "001001";
        when "0101111000100001" => data <= "001001";
        when "0101111000100010" => data <= "001001";
        when "0101111000100011" => data <= "001001";
        when "0101111000100100" => data <= "001001";
        when "0101111000100101" => data <= "001001";
        when "0101111000100110" => data <= "001001";
        when "0101111000100111" => data <= "001001";
        when "0101111000101000" => data <= "001001";
        when "0101111000101001" => data <= "001001";
        when "0101111000101010" => data <= "001001";
        when "0101111000101011" => data <= "001001";
        when "0101111000101100" => data <= "001001";
        when "0101111000101101" => data <= "001001";
        when "0101111000101110" => data <= "110000";
        when "0101111000101111" => data <= "110000";
        when "0101111001001010" => data <= "110000";
        when "0101111001011000" => data <= "110000";
        when "0101111001110001" => data <= "110000";
        when "0101111001110010" => data <= "001001";
        when "0101111001110011" => data <= "001001";
        when "0101111001110100" => data <= "001001";
        when "0101111001110101" => data <= "001001";
        when "0101111001110110" => data <= "001001";
        when "0101111001110111" => data <= "001001";
        when "0101111001111000" => data <= "001001";
        when "0101111001111001" => data <= "001001";
        when "0101111001111010" => data <= "001001";
        when "0101111001111011" => data <= "001001";
        when "0101111001111100" => data <= "001001";
        when "0101111001111101" => data <= "001001";
        when "0101111001111110" => data <= "001001";
        when "0101111001111111" => data <= "001001";
        when "0101111010000000" => data <= "001001";
        when "0101111010000001" => data <= "001001";
        when "0101111010000010" => data <= "001001";
        when "0101111010000011" => data <= "001001";
        when "0101111010000100" => data <= "001001";
        when "0101111010000101" => data <= "001001";
        when "0101111010000110" => data <= "001001";
        when "0101111010000111" => data <= "001001";
        when "0101111010001000" => data <= "110000";
        when "0101111010001001" => data <= "110000";
        when "0101111010011110" => data <= "110000";
        when "0101111010011111" => data <= "110000";
        when "0101111100000000" => data <= "110000";
        when "0101111100000001" => data <= "110000";
        when "0101111100011001" => data <= "110000";
        when "0101111100011010" => data <= "110000";
        when "0101111100011011" => data <= "001001";
        when "0101111100011100" => data <= "001001";
        when "0101111100011101" => data <= "001001";
        when "0101111100011110" => data <= "001001";
        when "0101111100011111" => data <= "001001";
        when "0101111100100000" => data <= "001001";
        when "0101111100100001" => data <= "001001";
        when "0101111100100010" => data <= "001001";
        when "0101111100100011" => data <= "001001";
        when "0101111100100100" => data <= "001001";
        when "0101111100100101" => data <= "001001";
        when "0101111100100110" => data <= "001001";
        when "0101111100100111" => data <= "001001";
        when "0101111100101000" => data <= "001001";
        when "0101111100101001" => data <= "001001";
        when "0101111100101010" => data <= "001001";
        when "0101111100101011" => data <= "001001";
        when "0101111100101100" => data <= "001001";
        when "0101111100101101" => data <= "001001";
        when "0101111100101110" => data <= "001001";
        when "0101111100101111" => data <= "001001";
        when "0101111100110000" => data <= "110000";
        when "0101111101001010" => data <= "110000";
        when "0101111101011000" => data <= "110000";
        when "0101111101101111" => data <= "110000";
        when "0101111101110000" => data <= "110000";
        when "0101111101110001" => data <= "001001";
        when "0101111101110010" => data <= "001001";
        when "0101111101110011" => data <= "001001";
        when "0101111101110100" => data <= "001001";
        when "0101111101110101" => data <= "001001";
        when "0101111101110110" => data <= "001001";
        when "0101111101110111" => data <= "001001";
        when "0101111101111000" => data <= "001001";
        when "0101111101111001" => data <= "001001";
        when "0101111101111010" => data <= "001001";
        when "0101111101111011" => data <= "001001";
        when "0101111101111100" => data <= "001001";
        when "0101111101111101" => data <= "001001";
        when "0101111101111110" => data <= "001001";
        when "0101111101111111" => data <= "001001";
        when "0101111110000000" => data <= "001001";
        when "0101111110000001" => data <= "001001";
        when "0101111110000010" => data <= "001001";
        when "0101111110000011" => data <= "001001";
        when "0101111110000100" => data <= "001001";
        when "0101111110000101" => data <= "110000";
        when "0101111110000110" => data <= "110000";
        when "0101111110000111" => data <= "110000";
        when "0101111110011110" => data <= "110000";
        when "0101111110011111" => data <= "110000";
        when "0110000000000000" => data <= "110000";
        when "0110000000000001" => data <= "110000";
        when "0110000000001000" => data <= "111111";
        when "0110000000001100" => data <= "111111";
        when "0110000000010000" => data <= "111111";
        when "0110000000011011" => data <= "110000";
        when "0110000000011100" => data <= "110000";
        when "0110000000011101" => data <= "001001";
        when "0110000000011110" => data <= "001001";
        when "0110000000011111" => data <= "001001";
        when "0110000000100000" => data <= "001001";
        when "0110000000100001" => data <= "001001";
        when "0110000000100010" => data <= "001001";
        when "0110000000100011" => data <= "001001";
        when "0110000000100100" => data <= "001001";
        when "0110000000100101" => data <= "001001";
        when "0110000000100110" => data <= "001001";
        when "0110000000100111" => data <= "001001";
        when "0110000000101000" => data <= "001001";
        when "0110000000101001" => data <= "001001";
        when "0110000000101010" => data <= "001001";
        when "0110000000101011" => data <= "001001";
        when "0110000000101100" => data <= "001001";
        when "0110000000101101" => data <= "001001";
        when "0110000000101110" => data <= "001001";
        when "0110000000101111" => data <= "001001";
        when "0110000000110000" => data <= "001001";
        when "0110000000110001" => data <= "110000";
        when "0110000001001010" => data <= "110000";
        when "0110000001011000" => data <= "110000";
        when "0110000001101110" => data <= "110000";
        when "0110000001101111" => data <= "001001";
        when "0110000001110000" => data <= "001001";
        when "0110000001110001" => data <= "001001";
        when "0110000001110010" => data <= "001001";
        when "0110000001110011" => data <= "001001";
        when "0110000001110100" => data <= "001001";
        when "0110000001110101" => data <= "001001";
        when "0110000001110110" => data <= "001001";
        when "0110000001110111" => data <= "001001";
        when "0110000001111000" => data <= "001001";
        when "0110000001111001" => data <= "001001";
        when "0110000001111010" => data <= "001001";
        when "0110000001111011" => data <= "001001";
        when "0110000001111100" => data <= "001001";
        when "0110000001111101" => data <= "001001";
        when "0110000001111110" => data <= "001001";
        when "0110000001111111" => data <= "001001";
        when "0110000010000000" => data <= "001001";
        when "0110000010000001" => data <= "001001";
        when "0110000010000010" => data <= "001001";
        when "0110000010000011" => data <= "110000";
        when "0110000010000100" => data <= "110000";
        when "0110000010001111" => data <= "111111";
        when "0110000010010011" => data <= "111111";
        when "0110000010010111" => data <= "111111";
        when "0110000010011110" => data <= "110000";
        when "0110000010011111" => data <= "110000";
        when "0110000100000000" => data <= "110000";
        when "0110000100000001" => data <= "110000";
        when "0110000100001001" => data <= "111111";
        when "0110000100001100" => data <= "111111";
        when "0110000100001111" => data <= "111111";
        when "0110000100011101" => data <= "110000";
        when "0110000100011110" => data <= "110000";
        when "0110000100011111" => data <= "001001";
        when "0110000100100000" => data <= "001001";
        when "0110000100100001" => data <= "001001";
        when "0110000100100010" => data <= "001001";
        when "0110000100100011" => data <= "001001";
        when "0110000100100100" => data <= "001001";
        when "0110000100100101" => data <= "001001";
        when "0110000100100110" => data <= "001001";
        when "0110000100100111" => data <= "001001";
        when "0110000100101000" => data <= "001001";
        when "0110000100101001" => data <= "001001";
        when "0110000100101010" => data <= "001001";
        when "0110000100101011" => data <= "001001";
        when "0110000100101100" => data <= "001001";
        when "0110000100101101" => data <= "001001";
        when "0110000100101110" => data <= "001001";
        when "0110000100101111" => data <= "001001";
        when "0110000100110000" => data <= "001001";
        when "0110000100110001" => data <= "001001";
        when "0110000100110010" => data <= "110000";
        when "0110000100110011" => data <= "110000";
        when "0110000101001010" => data <= "110000";
        when "0110000101011000" => data <= "110000";
        when "0110000101101101" => data <= "110000";
        when "0110000101101110" => data <= "001001";
        when "0110000101101111" => data <= "001001";
        when "0110000101110000" => data <= "001001";
        when "0110000101110001" => data <= "001001";
        when "0110000101110010" => data <= "001001";
        when "0110000101110011" => data <= "001001";
        when "0110000101110100" => data <= "001001";
        when "0110000101110101" => data <= "001001";
        when "0110000101110110" => data <= "001001";
        when "0110000101110111" => data <= "001001";
        when "0110000101111000" => data <= "001001";
        when "0110000101111001" => data <= "001001";
        when "0110000101111010" => data <= "001001";
        when "0110000101111011" => data <= "001001";
        when "0110000101111100" => data <= "001001";
        when "0110000101111101" => data <= "001001";
        when "0110000101111110" => data <= "001001";
        when "0110000101111111" => data <= "001001";
        when "0110000110000000" => data <= "001001";
        when "0110000110000001" => data <= "110000";
        when "0110000110000010" => data <= "110000";
        when "0110000110010000" => data <= "111111";
        when "0110000110010011" => data <= "111111";
        when "0110000110010110" => data <= "111111";
        when "0110000110011110" => data <= "110000";
        when "0110000110011111" => data <= "110000";
        when "0110001000000000" => data <= "110000";
        when "0110001000000001" => data <= "110000";
        when "0110001000001010" => data <= "111111";
        when "0110001000001100" => data <= "111111";
        when "0110001000001110" => data <= "111111";
        when "0110001000011111" => data <= "110000";
        when "0110001000100000" => data <= "110000";
        when "0110001000100001" => data <= "110000";
        when "0110001000100010" => data <= "001001";
        when "0110001000100011" => data <= "001001";
        when "0110001000100100" => data <= "001001";
        when "0110001000100101" => data <= "001001";
        when "0110001000100110" => data <= "001001";
        when "0110001000100111" => data <= "001001";
        when "0110001000101000" => data <= "001001";
        when "0110001000101001" => data <= "001001";
        when "0110001000101010" => data <= "001001";
        when "0110001000101011" => data <= "001001";
        when "0110001000101100" => data <= "001001";
        when "0110001000101101" => data <= "001001";
        when "0110001000101110" => data <= "001001";
        when "0110001000101111" => data <= "001001";
        when "0110001000110000" => data <= "001001";
        when "0110001000110001" => data <= "001001";
        when "0110001000110010" => data <= "001001";
        when "0110001000110011" => data <= "001001";
        when "0110001000110100" => data <= "110000";
        when "0110001001001010" => data <= "110000";
        when "0110001001010101" => data <= "110000";
        when "0110001001010110" => data <= "110000";
        when "0110001001010111" => data <= "110000";
        when "0110001001011000" => data <= "110000";
        when "0110001001101100" => data <= "110000";
        when "0110001001101101" => data <= "001001";
        when "0110001001101110" => data <= "001001";
        when "0110001001101111" => data <= "001001";
        when "0110001001110000" => data <= "001001";
        when "0110001001110001" => data <= "001001";
        when "0110001001110010" => data <= "001001";
        when "0110001001110011" => data <= "001001";
        when "0110001001110100" => data <= "001001";
        when "0110001001110101" => data <= "001001";
        when "0110001001110110" => data <= "001001";
        when "0110001001110111" => data <= "001001";
        when "0110001001111000" => data <= "001001";
        when "0110001001111001" => data <= "001001";
        when "0110001001111010" => data <= "001001";
        when "0110001001111011" => data <= "001001";
        when "0110001001111100" => data <= "001001";
        when "0110001001111101" => data <= "001001";
        when "0110001001111110" => data <= "001001";
        when "0110001001111111" => data <= "110000";
        when "0110001010000000" => data <= "110000";
        when "0110001010010001" => data <= "111111";
        when "0110001010010011" => data <= "111111";
        when "0110001010010101" => data <= "111111";
        when "0110001010011110" => data <= "110000";
        when "0110001010011111" => data <= "110000";
        when "0110001100000000" => data <= "110000";
        when "0110001100000001" => data <= "110000";
        when "0110001100001000" => data <= "111111";
        when "0110001100001011" => data <= "111111";
        when "0110001100001100" => data <= "111111";
        when "0110001100001101" => data <= "111111";
        when "0110001100010000" => data <= "111111";
        when "0110001100100010" => data <= "110000";
        when "0110001100100011" => data <= "110000";
        when "0110001100100100" => data <= "001001";
        when "0110001100100101" => data <= "001001";
        when "0110001100100110" => data <= "001001";
        when "0110001100100111" => data <= "001001";
        when "0110001100101000" => data <= "001001";
        when "0110001100101001" => data <= "001001";
        when "0110001100101010" => data <= "001001";
        when "0110001100101011" => data <= "001001";
        when "0110001100101100" => data <= "001001";
        when "0110001100101101" => data <= "001001";
        when "0110001100101110" => data <= "001001";
        when "0110001100101111" => data <= "001001";
        when "0110001100110000" => data <= "001001";
        when "0110001100110001" => data <= "001001";
        when "0110001100110010" => data <= "001001";
        when "0110001100110011" => data <= "001001";
        when "0110001100110100" => data <= "001001";
        when "0110001100110101" => data <= "110000";
        when "0110001101001010" => data <= "110000";
        when "0110001101010101" => data <= "110000";
        when "0110001101011000" => data <= "110000";
        when "0110001101101010" => data <= "110000";
        when "0110001101101011" => data <= "110000";
        when "0110001101101100" => data <= "001001";
        when "0110001101101101" => data <= "001001";
        when "0110001101101110" => data <= "001001";
        when "0110001101101111" => data <= "001001";
        when "0110001101110000" => data <= "001001";
        when "0110001101110001" => data <= "001001";
        when "0110001101110010" => data <= "001001";
        when "0110001101110011" => data <= "001001";
        when "0110001101110100" => data <= "001001";
        when "0110001101110101" => data <= "001001";
        when "0110001101110110" => data <= "001001";
        when "0110001101110111" => data <= "001001";
        when "0110001101111000" => data <= "001001";
        when "0110001101111001" => data <= "001001";
        when "0110001101111010" => data <= "001001";
        when "0110001101111011" => data <= "001001";
        when "0110001101111100" => data <= "001001";
        when "0110001101111101" => data <= "110000";
        when "0110001101111110" => data <= "110000";
        when "0110001110001111" => data <= "111111";
        when "0110001110010010" => data <= "111111";
        when "0110001110010011" => data <= "111111";
        when "0110001110010100" => data <= "111111";
        when "0110001110010111" => data <= "111111";
        when "0110001110011110" => data <= "110000";
        when "0110001110011111" => data <= "110000";
        when "0110010000000000" => data <= "110000";
        when "0110010000000001" => data <= "110000";
        when "0110010000000110" => data <= "111111";
        when "0110010000001000" => data <= "111111";
        when "0110010000001100" => data <= "111111";
        when "0110010000010000" => data <= "111111";
        when "0110010000010010" => data <= "111111";
        when "0110010000100100" => data <= "110000";
        when "0110010000100101" => data <= "110000";
        when "0110010000100110" => data <= "001001";
        when "0110010000100111" => data <= "001001";
        when "0110010000101000" => data <= "001001";
        when "0110010000101001" => data <= "001001";
        when "0110010000101010" => data <= "001001";
        when "0110010000101011" => data <= "001001";
        when "0110010000101100" => data <= "001001";
        when "0110010000101101" => data <= "001001";
        when "0110010000101110" => data <= "001001";
        when "0110010000101111" => data <= "001001";
        when "0110010000110000" => data <= "001001";
        when "0110010000110001" => data <= "001001";
        when "0110010000110010" => data <= "001001";
        when "0110010000110011" => data <= "001001";
        when "0110010000110100" => data <= "001001";
        when "0110010000110101" => data <= "001001";
        when "0110010000110110" => data <= "110000";
        when "0110010000110111" => data <= "110000";
        when "0110010001000110" => data <= "110000";
        when "0110010001000111" => data <= "110000";
        when "0110010001001000" => data <= "110000";
        when "0110010001001001" => data <= "110000";
        when "0110010001001010" => data <= "110000";
        when "0110010001010101" => data <= "110000";
        when "0110010001011000" => data <= "110000";
        when "0110010001101001" => data <= "110000";
        when "0110010001101010" => data <= "001001";
        when "0110010001101011" => data <= "001001";
        when "0110010001101100" => data <= "001001";
        when "0110010001101101" => data <= "001001";
        when "0110010001101110" => data <= "001001";
        when "0110010001101111" => data <= "001001";
        when "0110010001110000" => data <= "001001";
        when "0110010001110001" => data <= "001001";
        when "0110010001110010" => data <= "001001";
        when "0110010001110011" => data <= "001001";
        when "0110010001110100" => data <= "001001";
        when "0110010001110101" => data <= "001001";
        when "0110010001110110" => data <= "001001";
        when "0110010001110111" => data <= "001001";
        when "0110010001111000" => data <= "001001";
        when "0110010001111001" => data <= "001001";
        when "0110010001111010" => data <= "110000";
        when "0110010001111011" => data <= "110000";
        when "0110010001111100" => data <= "110000";
        when "0110010010001101" => data <= "111111";
        when "0110010010001111" => data <= "111111";
        when "0110010010010011" => data <= "111111";
        when "0110010010010111" => data <= "111111";
        when "0110010010011001" => data <= "111111";
        when "0110010010011110" => data <= "110000";
        when "0110010010011111" => data <= "110000";
        when "0110010100000000" => data <= "110000";
        when "0110010100000001" => data <= "110000";
        when "0110010100000111" => data <= "111111";
        when "0110010100001000" => data <= "111111";
        when "0110010100001100" => data <= "111111";
        when "0110010100010000" => data <= "111111";
        when "0110010100010001" => data <= "111111";
        when "0110010100100110" => data <= "110000";
        when "0110010100100111" => data <= "110000";
        when "0110010100101000" => data <= "001001";
        when "0110010100101001" => data <= "001001";
        when "0110010100101010" => data <= "001001";
        when "0110010100101011" => data <= "001001";
        when "0110010100101100" => data <= "001001";
        when "0110010100101101" => data <= "001001";
        when "0110010100101110" => data <= "001001";
        when "0110010100101111" => data <= "001001";
        when "0110010100110000" => data <= "001001";
        when "0110010100110001" => data <= "001001";
        when "0110010100110010" => data <= "001001";
        when "0110010100110011" => data <= "001001";
        when "0110010100110100" => data <= "001001";
        when "0110010100110101" => data <= "001001";
        when "0110010100110110" => data <= "001001";
        when "0110010100110111" => data <= "001001";
        when "0110010100111000" => data <= "110000";
        when "0110010101000110" => data <= "110000";
        when "0110010101001001" => data <= "110000";
        when "0110010101001010" => data <= "110000";
        when "0110010101010100" => data <= "110000";
        when "0110010101011000" => data <= "110000";
        when "0110010101101000" => data <= "110000";
        when "0110010101101001" => data <= "001001";
        when "0110010101101010" => data <= "001001";
        when "0110010101101011" => data <= "001001";
        when "0110010101101100" => data <= "001001";
        when "0110010101101101" => data <= "001001";
        when "0110010101101110" => data <= "001001";
        when "0110010101101111" => data <= "001001";
        when "0110010101110000" => data <= "001001";
        when "0110010101110001" => data <= "001001";
        when "0110010101110010" => data <= "001001";
        when "0110010101110011" => data <= "001001";
        when "0110010101110100" => data <= "001001";
        when "0110010101110101" => data <= "001001";
        when "0110010101110110" => data <= "001001";
        when "0110010101110111" => data <= "001001";
        when "0110010101111000" => data <= "110000";
        when "0110010101111001" => data <= "110000";
        when "0110010110001110" => data <= "111111";
        when "0110010110001111" => data <= "111111";
        when "0110010110010011" => data <= "111111";
        when "0110010110010111" => data <= "111111";
        when "0110010110011000" => data <= "111111";
        when "0110010110011110" => data <= "110000";
        when "0110010110011111" => data <= "110000";
        when "0110011000000000" => data <= "110000";
        when "0110011000000001" => data <= "110000";
        when "0110011000000100" => data <= "111111";
        when "0110011000000101" => data <= "111111";
        when "0110011000000110" => data <= "111111";
        when "0110011000000111" => data <= "111111";
        when "0110011000001000" => data <= "111111";
        when "0110011000001100" => data <= "111111";
        when "0110011000010000" => data <= "111111";
        when "0110011000010001" => data <= "111111";
        when "0110011000010010" => data <= "111111";
        when "0110011000010011" => data <= "111111";
        when "0110011000010100" => data <= "111111";
        when "0110011000101000" => data <= "110000";
        when "0110011000101001" => data <= "110000";
        when "0110011000101010" => data <= "110000";
        when "0110011000101011" => data <= "001001";
        when "0110011000101100" => data <= "001001";
        when "0110011000101101" => data <= "001001";
        when "0110011000101110" => data <= "001001";
        when "0110011000101111" => data <= "001001";
        when "0110011000110000" => data <= "001001";
        when "0110011000110001" => data <= "001001";
        when "0110011000110010" => data <= "001001";
        when "0110011000110011" => data <= "001001";
        when "0110011000110100" => data <= "001001";
        when "0110011000110101" => data <= "001001";
        when "0110011000110110" => data <= "001001";
        when "0110011000110111" => data <= "001001";
        when "0110011000111000" => data <= "001001";
        when "0110011000111001" => data <= "110000";
        when "0110011001000101" => data <= "110000";
        when "0110011001000110" => data <= "110000";
        when "0110011001001001" => data <= "110000";
        when "0110011001001010" => data <= "110000";
        when "0110011001010100" => data <= "110000";
        when "0110011001011000" => data <= "110000";
        when "0110011001100110" => data <= "110000";
        when "0110011001100111" => data <= "110000";
        when "0110011001101000" => data <= "001001";
        when "0110011001101001" => data <= "001001";
        when "0110011001101010" => data <= "001001";
        when "0110011001101011" => data <= "001001";
        when "0110011001101100" => data <= "001001";
        when "0110011001101101" => data <= "001001";
        when "0110011001101110" => data <= "001001";
        when "0110011001101111" => data <= "001001";
        when "0110011001110000" => data <= "001001";
        when "0110011001110001" => data <= "001001";
        when "0110011001110010" => data <= "001001";
        when "0110011001110011" => data <= "001001";
        when "0110011001110100" => data <= "001001";
        when "0110011001110101" => data <= "001001";
        when "0110011001110110" => data <= "110000";
        when "0110011001110111" => data <= "110000";
        when "0110011010001011" => data <= "111111";
        when "0110011010001100" => data <= "111111";
        when "0110011010001101" => data <= "111111";
        when "0110011010001110" => data <= "111111";
        when "0110011010001111" => data <= "111111";
        when "0110011010010011" => data <= "111111";
        when "0110011010010111" => data <= "111111";
        when "0110011010011000" => data <= "111111";
        when "0110011010011001" => data <= "111111";
        when "0110011010011010" => data <= "111111";
        when "0110011010011011" => data <= "111111";
        when "0110011010011110" => data <= "110000";
        when "0110011010011111" => data <= "110000";
        when "0110011100000000" => data <= "110000";
        when "0110011100000001" => data <= "110000";
        when "0110011100001001" => data <= "111111";
        when "0110011100001100" => data <= "111111";
        when "0110011100001111" => data <= "111111";
        when "0110011100101011" => data <= "110000";
        when "0110011100101100" => data <= "110000";
        when "0110011100101101" => data <= "001001";
        when "0110011100101110" => data <= "001001";
        when "0110011100101111" => data <= "001001";
        when "0110011100110000" => data <= "001001";
        when "0110011100110001" => data <= "001001";
        when "0110011100110010" => data <= "001001";
        when "0110011100110011" => data <= "001001";
        when "0110011100110100" => data <= "001001";
        when "0110011100110101" => data <= "001001";
        when "0110011100110110" => data <= "001001";
        when "0110011100110111" => data <= "001001";
        when "0110011100111000" => data <= "001001";
        when "0110011100111001" => data <= "001001";
        when "0110011100111010" => data <= "110000";
        when "0110011100111011" => data <= "110000";
        when "0110011101000101" => data <= "110000";
        when "0110011101001010" => data <= "110000";
        when "0110011101010100" => data <= "110000";
        when "0110011101011000" => data <= "110000";
        when "0110011101100101" => data <= "110000";
        when "0110011101100110" => data <= "001001";
        when "0110011101100111" => data <= "001001";
        when "0110011101101000" => data <= "001001";
        when "0110011101101001" => data <= "001001";
        when "0110011101101010" => data <= "001001";
        when "0110011101101011" => data <= "001001";
        when "0110011101101100" => data <= "001001";
        when "0110011101101101" => data <= "001001";
        when "0110011101101110" => data <= "001001";
        when "0110011101101111" => data <= "001001";
        when "0110011101110000" => data <= "001001";
        when "0110011101110001" => data <= "001001";
        when "0110011101110010" => data <= "001001";
        when "0110011101110011" => data <= "001001";
        when "0110011101110100" => data <= "110000";
        when "0110011101110101" => data <= "110000";
        when "0110011110010000" => data <= "111111";
        when "0110011110010011" => data <= "111111";
        when "0110011110010110" => data <= "111111";
        when "0110011110011110" => data <= "110000";
        when "0110011110011111" => data <= "110000";
        when "0110100000000000" => data <= "110000";
        when "0110100000000001" => data <= "110000";
        when "0110100000000101" => data <= "111111";
        when "0110100000001010" => data <= "111111";
        when "0110100000001100" => data <= "111111";
        when "0110100000001110" => data <= "111111";
        when "0110100000010011" => data <= "111111";
        when "0110100000101101" => data <= "110000";
        when "0110100000101110" => data <= "110000";
        when "0110100000101111" => data <= "001001";
        when "0110100000110000" => data <= "001001";
        when "0110100000110001" => data <= "001001";
        when "0110100000110010" => data <= "001001";
        when "0110100000110011" => data <= "001001";
        when "0110100000110100" => data <= "001001";
        when "0110100000110101" => data <= "001001";
        when "0110100000110110" => data <= "001001";
        when "0110100000110111" => data <= "001001";
        when "0110100000111000" => data <= "001001";
        when "0110100000111001" => data <= "001001";
        when "0110100000111010" => data <= "001001";
        when "0110100000111011" => data <= "001001";
        when "0110100000111100" => data <= "110000";
        when "0110100001000101" => data <= "110000";
        when "0110100001001010" => data <= "110000";
        when "0110100001010100" => data <= "110000";
        when "0110100001011000" => data <= "110000";
        when "0110100001100100" => data <= "110000";
        when "0110100001100101" => data <= "001001";
        when "0110100001100110" => data <= "001001";
        when "0110100001100111" => data <= "001001";
        when "0110100001101000" => data <= "001001";
        when "0110100001101001" => data <= "001001";
        when "0110100001101010" => data <= "001001";
        when "0110100001101011" => data <= "001001";
        when "0110100001101100" => data <= "001001";
        when "0110100001101101" => data <= "001001";
        when "0110100001101110" => data <= "001001";
        when "0110100001101111" => data <= "001001";
        when "0110100001110000" => data <= "001001";
        when "0110100001110001" => data <= "110000";
        when "0110100001110010" => data <= "110000";
        when "0110100001110011" => data <= "110000";
        when "0110100010001100" => data <= "111111";
        when "0110100010010001" => data <= "111111";
        when "0110100010010011" => data <= "111111";
        when "0110100010010101" => data <= "111111";
        when "0110100010011010" => data <= "111111";
        when "0110100010011110" => data <= "110000";
        when "0110100010011111" => data <= "110000";
        when "0110100100000000" => data <= "110000";
        when "0110100100000001" => data <= "110000";
        when "0110100100000110" => data <= "111111";
        when "0110100100001011" => data <= "111111";
        when "0110100100001100" => data <= "111111";
        when "0110100100001101" => data <= "111111";
        when "0110100100010010" => data <= "111111";
        when "0110100100101111" => data <= "110000";
        when "0110100100110000" => data <= "110000";
        when "0110100100110001" => data <= "001001";
        when "0110100100110010" => data <= "001001";
        when "0110100100110011" => data <= "001001";
        when "0110100100110100" => data <= "001001";
        when "0110100100110101" => data <= "001001";
        when "0110100100110110" => data <= "001001";
        when "0110100100110111" => data <= "001001";
        when "0110100100111000" => data <= "001001";
        when "0110100100111001" => data <= "001001";
        when "0110100100111010" => data <= "001001";
        when "0110100100111011" => data <= "001001";
        when "0110100100111100" => data <= "001001";
        when "0110100100111101" => data <= "110000";
        when "0110100101000101" => data <= "110000";
        when "0110100101000110" => data <= "110000";
        when "0110100101001010" => data <= "110000";
        when "0110100101010100" => data <= "110000";
        when "0110100101010110" => data <= "110000";
        when "0110100101010111" => data <= "110000";
        when "0110100101011000" => data <= "110000";
        when "0110100101100010" => data <= "110000";
        when "0110100101100011" => data <= "110000";
        when "0110100101100100" => data <= "001001";
        when "0110100101100101" => data <= "001001";
        when "0110100101100110" => data <= "001001";
        when "0110100101100111" => data <= "001001";
        when "0110100101101000" => data <= "001001";
        when "0110100101101001" => data <= "001001";
        when "0110100101101010" => data <= "001001";
        when "0110100101101011" => data <= "001001";
        when "0110100101101100" => data <= "001001";
        when "0110100101101101" => data <= "001001";
        when "0110100101101110" => data <= "001001";
        when "0110100101101111" => data <= "110000";
        when "0110100101110000" => data <= "110000";
        when "0110100110001101" => data <= "111111";
        when "0110100110010010" => data <= "111111";
        when "0110100110010011" => data <= "111111";
        when "0110100110010100" => data <= "111111";
        when "0110100110011001" => data <= "111111";
        when "0110100110011110" => data <= "110000";
        when "0110100110011111" => data <= "110000";
        when "0110101000000000" => data <= "110000";
        when "0110101000000001" => data <= "110000";
        when "0110101000000011" => data <= "111111";
        when "0110101000000100" => data <= "111111";
        when "0110101000000101" => data <= "111111";
        when "0110101000000110" => data <= "111111";
        when "0110101000000111" => data <= "111111";
        when "0110101000001000" => data <= "111111";
        when "0110101000001001" => data <= "111111";
        when "0110101000001010" => data <= "111111";
        when "0110101000001011" => data <= "111111";
        when "0110101000001100" => data <= "111111";
        when "0110101000001101" => data <= "111111";
        when "0110101000001110" => data <= "111111";
        when "0110101000001111" => data <= "111111";
        when "0110101000010000" => data <= "111111";
        when "0110101000010001" => data <= "111111";
        when "0110101000010010" => data <= "111111";
        when "0110101000010011" => data <= "111111";
        when "0110101000010100" => data <= "111111";
        when "0110101000010101" => data <= "111111";
        when "0110101000110001" => data <= "110000";
        when "0110101000110010" => data <= "110000";
        when "0110101000110011" => data <= "110000";
        when "0110101000110100" => data <= "001001";
        when "0110101000110101" => data <= "001001";
        when "0110101000110110" => data <= "001001";
        when "0110101000110111" => data <= "001001";
        when "0110101000111000" => data <= "001001";
        when "0110101000111001" => data <= "001001";
        when "0110101000111010" => data <= "001001";
        when "0110101000111011" => data <= "001001";
        when "0110101000111100" => data <= "001001";
        when "0110101000111101" => data <= "001001";
        when "0110101000111110" => data <= "110000";
        when "0110101000111111" => data <= "110000";
        when "0110101001000110" => data <= "110000";
        when "0110101001001010" => data <= "110000";
        when "0110101001010100" => data <= "110000";
        when "0110101001010101" => data <= "110000";
        when "0110101001010110" => data <= "110000";
        when "0110101001100001" => data <= "110000";
        when "0110101001100010" => data <= "001001";
        when "0110101001100011" => data <= "001001";
        when "0110101001100100" => data <= "001001";
        when "0110101001100101" => data <= "001001";
        when "0110101001100110" => data <= "001001";
        when "0110101001100111" => data <= "001001";
        when "0110101001101000" => data <= "001001";
        when "0110101001101001" => data <= "001001";
        when "0110101001101010" => data <= "001001";
        when "0110101001101011" => data <= "001001";
        when "0110101001101100" => data <= "001001";
        when "0110101001101101" => data <= "110000";
        when "0110101001101110" => data <= "110000";
        when "0110101010001010" => data <= "111111";
        when "0110101010001011" => data <= "111111";
        when "0110101010001100" => data <= "111111";
        when "0110101010001101" => data <= "111111";
        when "0110101010001110" => data <= "111111";
        when "0110101010001111" => data <= "111111";
        when "0110101010010000" => data <= "111111";
        when "0110101010010001" => data <= "111111";
        when "0110101010010010" => data <= "111111";
        when "0110101010010011" => data <= "111111";
        when "0110101010010100" => data <= "111111";
        when "0110101010010101" => data <= "111111";
        when "0110101010010110" => data <= "111111";
        when "0110101010010111" => data <= "111111";
        when "0110101010011000" => data <= "111111";
        when "0110101010011001" => data <= "111111";
        when "0110101010011010" => data <= "111111";
        when "0110101010011011" => data <= "111111";
        when "0110101010011100" => data <= "111111";
        when "0110101010011110" => data <= "110000";
        when "0110101010011111" => data <= "110000";
        when "0110101100000000" => data <= "110000";
        when "0110101100000001" => data <= "110000";
        when "0110101100000110" => data <= "111111";
        when "0110101100001011" => data <= "111111";
        when "0110101100001100" => data <= "111111";
        when "0110101100001101" => data <= "111111";
        when "0110101100010010" => data <= "111111";
        when "0110101100110100" => data <= "110000";
        when "0110101100110101" => data <= "110000";
        when "0110101100110110" => data <= "001001";
        when "0110101100110111" => data <= "001001";
        when "0110101100111000" => data <= "001001";
        when "0110101100111001" => data <= "001001";
        when "0110101100111010" => data <= "001001";
        when "0110101100111011" => data <= "001001";
        when "0110101100111100" => data <= "001001";
        when "0110101100111101" => data <= "001001";
        when "0110101100111110" => data <= "001001";
        when "0110101100111111" => data <= "001001";
        when "0110101101000000" => data <= "110000";
        when "0110101101000110" => data <= "110000";
        when "0110101101000111" => data <= "110000";
        when "0110101101001010" => data <= "110000";
        when "0110101101100000" => data <= "110000";
        when "0110101101100001" => data <= "001001";
        when "0110101101100010" => data <= "001001";
        when "0110101101100011" => data <= "001001";
        when "0110101101100100" => data <= "001001";
        when "0110101101100101" => data <= "001001";
        when "0110101101100110" => data <= "001001";
        when "0110101101100111" => data <= "001001";
        when "0110101101101000" => data <= "001001";
        when "0110101101101001" => data <= "001001";
        when "0110101101101010" => data <= "001001";
        when "0110101101101011" => data <= "110000";
        when "0110101101101100" => data <= "110000";
        when "0110101110001101" => data <= "111111";
        when "0110101110010010" => data <= "111111";
        when "0110101110010011" => data <= "111111";
        when "0110101110010100" => data <= "111111";
        when "0110101110011001" => data <= "111111";
        when "0110101110011110" => data <= "110000";
        when "0110101110011111" => data <= "110000";
        when "0110110000000000" => data <= "110000";
        when "0110110000000001" => data <= "110000";
        when "0110110000000101" => data <= "111111";
        when "0110110000001010" => data <= "111111";
        when "0110110000001100" => data <= "111111";
        when "0110110000001110" => data <= "111111";
        when "0110110000010011" => data <= "111111";
        when "0110110000110110" => data <= "110000";
        when "0110110000110111" => data <= "110000";
        when "0110110000111000" => data <= "001001";
        when "0110110000111001" => data <= "001001";
        when "0110110000111010" => data <= "001001";
        when "0110110000111011" => data <= "001001";
        when "0110110000111100" => data <= "001001";
        when "0110110000111101" => data <= "001001";
        when "0110110000111110" => data <= "001001";
        when "0110110000111111" => data <= "001001";
        when "0110110001000000" => data <= "001001";
        when "0110110001000001" => data <= "110000";
        when "0110110001000111" => data <= "110000";
        when "0110110001001000" => data <= "110000";
        when "0110110001001001" => data <= "110000";
        when "0110110001001010" => data <= "110000";
        when "0110110001011110" => data <= "110000";
        when "0110110001011111" => data <= "110000";
        when "0110110001100000" => data <= "001001";
        when "0110110001100001" => data <= "001001";
        when "0110110001100010" => data <= "001001";
        when "0110110001100011" => data <= "001001";
        when "0110110001100100" => data <= "001001";
        when "0110110001100101" => data <= "001001";
        when "0110110001100110" => data <= "001001";
        when "0110110001100111" => data <= "001001";
        when "0110110001101000" => data <= "110000";
        when "0110110001101001" => data <= "110000";
        when "0110110001101010" => data <= "110000";
        when "0110110010001100" => data <= "111111";
        when "0110110010010001" => data <= "111111";
        when "0110110010010011" => data <= "111111";
        when "0110110010010101" => data <= "111111";
        when "0110110010011010" => data <= "111111";
        when "0110110010011110" => data <= "110000";
        when "0110110010011111" => data <= "110000";
        when "0110110100000000" => data <= "110000";
        when "0110110100000001" => data <= "110000";
        when "0110110100001001" => data <= "111111";
        when "0110110100001100" => data <= "111111";
        when "0110110100001111" => data <= "111111";
        when "0110110100111000" => data <= "110000";
        when "0110110100111001" => data <= "110000";
        when "0110110100111010" => data <= "001001";
        when "0110110100111011" => data <= "001001";
        when "0110110100111100" => data <= "001001";
        when "0110110100111101" => data <= "001001";
        when "0110110100111110" => data <= "001001";
        when "0110110100111111" => data <= "001001";
        when "0110110101000000" => data <= "001001";
        when "0110110101000001" => data <= "001001";
        when "0110110101000010" => data <= "110000";
        when "0110110101000011" => data <= "110000";
        when "0110110101011101" => data <= "110000";
        when "0110110101011110" => data <= "001001";
        when "0110110101011111" => data <= "001001";
        when "0110110101100000" => data <= "001001";
        when "0110110101100001" => data <= "001001";
        when "0110110101100010" => data <= "001001";
        when "0110110101100011" => data <= "001001";
        when "0110110101100100" => data <= "001001";
        when "0110110101100101" => data <= "001001";
        when "0110110101100110" => data <= "110000";
        when "0110110101100111" => data <= "110000";
        when "0110110110010000" => data <= "111111";
        when "0110110110010011" => data <= "111111";
        when "0110110110010110" => data <= "111111";
        when "0110110110011110" => data <= "110000";
        when "0110110110011111" => data <= "110000";
        when "0110111000000000" => data <= "110000";
        when "0110111000000001" => data <= "110000";
        when "0110111000000100" => data <= "111111";
        when "0110111000000101" => data <= "111111";
        when "0110111000000110" => data <= "111111";
        when "0110111000000111" => data <= "111111";
        when "0110111000001000" => data <= "111111";
        when "0110111000001100" => data <= "111111";
        when "0110111000010000" => data <= "111111";
        when "0110111000010001" => data <= "111111";
        when "0110111000010010" => data <= "111111";
        when "0110111000010011" => data <= "111111";
        when "0110111000010100" => data <= "111111";
        when "0110111000111010" => data <= "110000";
        when "0110111000111011" => data <= "110000";
        when "0110111000111100" => data <= "110000";
        when "0110111000111101" => data <= "001001";
        when "0110111000111110" => data <= "001001";
        when "0110111000111111" => data <= "001001";
        when "0110111001000000" => data <= "001001";
        when "0110111001000001" => data <= "001001";
        when "0110111001000010" => data <= "001001";
        when "0110111001000011" => data <= "001001";
        when "0110111001000100" => data <= "110000";
        when "0110111001011100" => data <= "110000";
        when "0110111001011101" => data <= "001001";
        when "0110111001011110" => data <= "001001";
        when "0110111001011111" => data <= "001001";
        when "0110111001100000" => data <= "001001";
        when "0110111001100001" => data <= "001001";
        when "0110111001100010" => data <= "001001";
        when "0110111001100011" => data <= "001001";
        when "0110111001100100" => data <= "110000";
        when "0110111001100101" => data <= "110000";
        when "0110111010001011" => data <= "111111";
        when "0110111010001100" => data <= "111111";
        when "0110111010001101" => data <= "111111";
        when "0110111010001110" => data <= "111111";
        when "0110111010001111" => data <= "111111";
        when "0110111010010011" => data <= "111111";
        when "0110111010010111" => data <= "111111";
        when "0110111010011000" => data <= "111111";
        when "0110111010011001" => data <= "111111";
        when "0110111010011010" => data <= "111111";
        when "0110111010011011" => data <= "111111";
        when "0110111010011110" => data <= "110000";
        when "0110111010011111" => data <= "110000";
        when "0110111100000000" => data <= "110000";
        when "0110111100000001" => data <= "110000";
        when "0110111100000111" => data <= "111111";
        when "0110111100001000" => data <= "111111";
        when "0110111100001100" => data <= "111111";
        when "0110111100010000" => data <= "111111";
        when "0110111100010001" => data <= "111111";
        when "0110111100111101" => data <= "110000";
        when "0110111100111110" => data <= "110000";
        when "0110111100111111" => data <= "001001";
        when "0110111101000000" => data <= "001001";
        when "0110111101000001" => data <= "001001";
        when "0110111101000010" => data <= "001001";
        when "0110111101000011" => data <= "001001";
        when "0110111101000100" => data <= "001001";
        when "0110111101000101" => data <= "110000";
        when "0110111101011010" => data <= "110000";
        when "0110111101011011" => data <= "110000";
        when "0110111101011100" => data <= "001001";
        when "0110111101011101" => data <= "001001";
        when "0110111101011110" => data <= "001001";
        when "0110111101011111" => data <= "001001";
        when "0110111101100000" => data <= "001001";
        when "0110111101100001" => data <= "001001";
        when "0110111101100010" => data <= "110000";
        when "0110111101100011" => data <= "110000";
        when "0110111110001110" => data <= "111111";
        when "0110111110001111" => data <= "111111";
        when "0110111110010011" => data <= "111111";
        when "0110111110010111" => data <= "111111";
        when "0110111110011000" => data <= "111111";
        when "0110111110011110" => data <= "110000";
        when "0110111110011111" => data <= "110000";
        when "0111000000000000" => data <= "110000";
        when "0111000000000001" => data <= "110000";
        when "0111000000000110" => data <= "111111";
        when "0111000000001000" => data <= "111111";
        when "0111000000001100" => data <= "111111";
        when "0111000000010000" => data <= "111111";
        when "0111000000010010" => data <= "111111";
        when "0111000000111111" => data <= "110000";
        when "0111000001000000" => data <= "110000";
        when "0111000001000001" => data <= "001001";
        when "0111000001000010" => data <= "001001";
        when "0111000001000011" => data <= "001001";
        when "0111000001000100" => data <= "001001";
        when "0111000001000101" => data <= "001001";
        when "0111000001000110" => data <= "110000";
        when "0111000001000111" => data <= "110000";
        when "0111000001011001" => data <= "110000";
        when "0111000001011010" => data <= "001001";
        when "0111000001011011" => data <= "001001";
        when "0111000001011100" => data <= "001001";
        when "0111000001011101" => data <= "001001";
        when "0111000001011110" => data <= "001001";
        when "0111000001011111" => data <= "001001";
        when "0111000001100000" => data <= "110000";
        when "0111000001100001" => data <= "110000";
        when "0111000010001101" => data <= "111111";
        when "0111000010001111" => data <= "111111";
        when "0111000010010011" => data <= "111111";
        when "0111000010010111" => data <= "111111";
        when "0111000010011001" => data <= "111111";
        when "0111000010011110" => data <= "110000";
        when "0111000010011111" => data <= "110000";
        when "0111000100000000" => data <= "110000";
        when "0111000100000001" => data <= "110000";
        when "0111000100001000" => data <= "111111";
        when "0111000100001011" => data <= "111111";
        when "0111000100001100" => data <= "111111";
        when "0111000100001101" => data <= "111111";
        when "0111000100010000" => data <= "111111";
        when "0111000101000001" => data <= "110000";
        when "0111000101000010" => data <= "110000";
        when "0111000101000011" => data <= "001001";
        when "0111000101000100" => data <= "001001";
        when "0111000101000101" => data <= "001001";
        when "0111000101000110" => data <= "001001";
        when "0111000101000111" => data <= "001001";
        when "0111000101001000" => data <= "110000";
        when "0111000101011000" => data <= "110000";
        when "0111000101011001" => data <= "001001";
        when "0111000101011010" => data <= "001001";
        when "0111000101011011" => data <= "001001";
        when "0111000101011100" => data <= "001001";
        when "0111000101011101" => data <= "110000";
        when "0111000101011110" => data <= "110000";
        when "0111000101011111" => data <= "110000";
        when "0111000110001111" => data <= "111111";
        when "0111000110010010" => data <= "111111";
        when "0111000110010011" => data <= "111111";
        when "0111000110010100" => data <= "111111";
        when "0111000110010111" => data <= "111111";
        when "0111000110011110" => data <= "110000";
        when "0111000110011111" => data <= "110000";
        when "0111001000000000" => data <= "110000";
        when "0111001000000001" => data <= "110000";
        when "0111001000001010" => data <= "111111";
        when "0111001000001100" => data <= "111111";
        when "0111001000001110" => data <= "111111";
        when "0111001001000011" => data <= "110000";
        when "0111001001000100" => data <= "110000";
        when "0111001001000101" => data <= "110000";
        when "0111001001000110" => data <= "001001";
        when "0111001001000111" => data <= "001001";
        when "0111001001001000" => data <= "001001";
        when "0111001001001001" => data <= "110000";
        when "0111001001010111" => data <= "110000";
        when "0111001001011000" => data <= "001001";
        when "0111001001011001" => data <= "001001";
        when "0111001001011010" => data <= "001001";
        when "0111001001011011" => data <= "110000";
        when "0111001001011100" => data <= "110000";
        when "0111001010010001" => data <= "111111";
        when "0111001010010011" => data <= "111111";
        when "0111001010010101" => data <= "111111";
        when "0111001010011110" => data <= "110000";
        when "0111001010011111" => data <= "110000";
        when "0111001100000000" => data <= "110000";
        when "0111001100000001" => data <= "110000";
        when "0111001100001001" => data <= "111111";
        when "0111001100001100" => data <= "111111";
        when "0111001100001111" => data <= "111111";
        when "0111001101000110" => data <= "110000";
        when "0111001101000111" => data <= "110000";
        when "0111001101001000" => data <= "001001";
        when "0111001101001001" => data <= "001001";
        when "0111001101001010" => data <= "110000";
        when "0111001101001011" => data <= "110000";
        when "0111001101010101" => data <= "110000";
        when "0111001101010110" => data <= "110000";
        when "0111001101010111" => data <= "001001";
        when "0111001101011000" => data <= "001001";
        when "0111001101011001" => data <= "110000";
        when "0111001101011010" => data <= "110000";
        when "0111001110010000" => data <= "111111";
        when "0111001110010011" => data <= "111111";
        when "0111001110010110" => data <= "111111";
        when "0111001110011110" => data <= "110000";
        when "0111001110011111" => data <= "110000";
        when "0111010000000000" => data <= "110000";
        when "0111010000000001" => data <= "110000";
        when "0111010000001000" => data <= "111111";
        when "0111010000001100" => data <= "111111";
        when "0111010000010000" => data <= "111111";
        when "0111010001001000" => data <= "110000";
        when "0111010001001001" => data <= "110000";
        when "0111010001001010" => data <= "001001";
        when "0111010001001011" => data <= "001001";
        when "0111010001001100" => data <= "110000";
        when "0111010001010100" => data <= "110000";
        when "0111010001010101" => data <= "001001";
        when "0111010001010110" => data <= "001001";
        when "0111010001010111" => data <= "110000";
        when "0111010001011000" => data <= "110000";
        when "0111010010001111" => data <= "111111";
        when "0111010010010011" => data <= "111111";
        when "0111010010010111" => data <= "111111";
        when "0111010010011110" => data <= "110000";
        when "0111010010011111" => data <= "110000";
        when "0111010100000000" => data <= "110000";
        when "0111010100000001" => data <= "110000";
        when "0111010101001010" => data <= "110000";
        when "0111010101001011" => data <= "110000";
        when "0111010101001100" => data <= "001001";
        when "0111010101001101" => data <= "110000";
        when "0111010101010011" => data <= "110000";
        when "0111010101010100" => data <= "110000";
        when "0111010101010101" => data <= "110000";
        when "0111010101010110" => data <= "110000";
        when "0111010110011110" => data <= "110000";
        when "0111010110011111" => data <= "110000";
        when "0111011000000000" => data <= "110000";
        when "0111011000000001" => data <= "110000";
        when "0111011000000010" => data <= "110000";
        when "0111011000000011" => data <= "110000";
        when "0111011000000100" => data <= "110000";
        when "0111011000000101" => data <= "110000";
        when "0111011000000110" => data <= "110000";
        when "0111011000000111" => data <= "110000";
        when "0111011000001000" => data <= "110000";
        when "0111011000001001" => data <= "110000";
        when "0111011000001010" => data <= "110000";
        when "0111011000001011" => data <= "110000";
        when "0111011000001100" => data <= "110000";
        when "0111011000001101" => data <= "110000";
        when "0111011000001110" => data <= "110000";
        when "0111011000001111" => data <= "110000";
        when "0111011000010000" => data <= "110000";
        when "0111011000010001" => data <= "110000";
        when "0111011000010010" => data <= "110000";
        when "0111011000010011" => data <= "110000";
        when "0111011000010100" => data <= "110000";
        when "0111011000010101" => data <= "110000";
        when "0111011000010110" => data <= "110000";
        when "0111011000010111" => data <= "110000";
        when "0111011000011000" => data <= "110000";
        when "0111011000011001" => data <= "110000";
        when "0111011000011010" => data <= "110000";
        when "0111011000011011" => data <= "110000";
        when "0111011000011100" => data <= "110000";
        when "0111011000011101" => data <= "110000";
        when "0111011000011110" => data <= "110000";
        when "0111011000011111" => data <= "110000";
        when "0111011000100000" => data <= "110000";
        when "0111011000100001" => data <= "110000";
        when "0111011000100010" => data <= "110000";
        when "0111011000100011" => data <= "110000";
        when "0111011000100100" => data <= "110000";
        when "0111011000100101" => data <= "110000";
        when "0111011000100110" => data <= "110000";
        when "0111011000100111" => data <= "110000";
        when "0111011000101000" => data <= "110000";
        when "0111011000101001" => data <= "110000";
        when "0111011000101010" => data <= "110000";
        when "0111011000101011" => data <= "110000";
        when "0111011000101100" => data <= "110000";
        when "0111011000101101" => data <= "110000";
        when "0111011000101110" => data <= "110000";
        when "0111011000101111" => data <= "110000";
        when "0111011000110000" => data <= "110000";
        when "0111011000110001" => data <= "110000";
        when "0111011000110010" => data <= "110000";
        when "0111011000110011" => data <= "110000";
        when "0111011000110100" => data <= "110000";
        when "0111011000110101" => data <= "110000";
        when "0111011000110110" => data <= "110000";
        when "0111011000110111" => data <= "110000";
        when "0111011000111000" => data <= "110000";
        when "0111011000111001" => data <= "110000";
        when "0111011000111010" => data <= "110000";
        when "0111011000111011" => data <= "110000";
        when "0111011000111100" => data <= "110000";
        when "0111011000111101" => data <= "110000";
        when "0111011000111110" => data <= "110000";
        when "0111011000111111" => data <= "110000";
        when "0111011001000000" => data <= "110000";
        when "0111011001000001" => data <= "110000";
        when "0111011001000010" => data <= "110000";
        when "0111011001000011" => data <= "110000";
        when "0111011001000100" => data <= "110000";
        when "0111011001000101" => data <= "110000";
        when "0111011001000110" => data <= "110000";
        when "0111011001000111" => data <= "110000";
        when "0111011001001000" => data <= "110000";
        when "0111011001001001" => data <= "110000";
        when "0111011001001010" => data <= "110000";
        when "0111011001001011" => data <= "110000";
        when "0111011001001100" => data <= "110000";
        when "0111011001001101" => data <= "110000";
        when "0111011001001110" => data <= "110000";
        when "0111011001001111" => data <= "110000";
        when "0111011001010000" => data <= "110000";
        when "0111011001010001" => data <= "110000";
        when "0111011001010010" => data <= "110000";
        when "0111011001010011" => data <= "110000";
        when "0111011001010100" => data <= "110000";
        when "0111011001010101" => data <= "110000";
        when "0111011001010110" => data <= "110000";
        when "0111011001010111" => data <= "110000";
        when "0111011001011000" => data <= "110000";
        when "0111011001011001" => data <= "110000";
        when "0111011001011010" => data <= "110000";
        when "0111011001011011" => data <= "110000";
        when "0111011001011100" => data <= "110000";
        when "0111011001011101" => data <= "110000";
        when "0111011001011110" => data <= "110000";
        when "0111011001011111" => data <= "110000";
        when "0111011001100000" => data <= "110000";
        when "0111011001100001" => data <= "110000";
        when "0111011001100010" => data <= "110000";
        when "0111011001100011" => data <= "110000";
        when "0111011001100100" => data <= "110000";
        when "0111011001100101" => data <= "110000";
        when "0111011001100110" => data <= "110000";
        when "0111011001100111" => data <= "110000";
        when "0111011001101000" => data <= "110000";
        when "0111011001101001" => data <= "110000";
        when "0111011001101010" => data <= "110000";
        when "0111011001101011" => data <= "110000";
        when "0111011001101100" => data <= "110000";
        when "0111011001101101" => data <= "110000";
        when "0111011001101110" => data <= "110000";
        when "0111011001101111" => data <= "110000";
        when "0111011001110000" => data <= "110000";
        when "0111011001110001" => data <= "110000";
        when "0111011001110010" => data <= "110000";
        when "0111011001110011" => data <= "110000";
        when "0111011001110100" => data <= "110000";
        when "0111011001110101" => data <= "110000";
        when "0111011001110110" => data <= "110000";
        when "0111011001110111" => data <= "110000";
        when "0111011001111000" => data <= "110000";
        when "0111011001111001" => data <= "110000";
        when "0111011001111010" => data <= "110000";
        when "0111011001111011" => data <= "110000";
        when "0111011001111100" => data <= "110000";
        when "0111011001111101" => data <= "110000";
        when "0111011001111110" => data <= "110000";
        when "0111011001111111" => data <= "110000";
        when "0111011010000000" => data <= "110000";
        when "0111011010000001" => data <= "110000";
        when "0111011010000010" => data <= "110000";
        when "0111011010000011" => data <= "110000";
        when "0111011010000100" => data <= "110000";
        when "0111011010000101" => data <= "110000";
        when "0111011010000110" => data <= "110000";
        when "0111011010000111" => data <= "110000";
        when "0111011010001000" => data <= "110000";
        when "0111011010001001" => data <= "110000";
        when "0111011010001010" => data <= "110000";
        when "0111011010001011" => data <= "110000";
        when "0111011010001100" => data <= "110000";
        when "0111011010001101" => data <= "110000";
        when "0111011010001110" => data <= "110000";
        when "0111011010001111" => data <= "110000";
        when "0111011010010000" => data <= "110000";
        when "0111011010010001" => data <= "110000";
        when "0111011010010010" => data <= "110000";
        when "0111011010010011" => data <= "110000";
        when "0111011010010100" => data <= "110000";
        when "0111011010010101" => data <= "110000";
        when "0111011010010110" => data <= "110000";
        when "0111011010010111" => data <= "110000";
        when "0111011010011000" => data <= "110000";
        when "0111011010011001" => data <= "110000";
        when "0111011010011010" => data <= "110000";
        when "0111011010011011" => data <= "110000";
        when "0111011010011100" => data <= "110000";
        when "0111011010011101" => data <= "110000";
        when "0111011010011110" => data <= "110000";
        when "0111011010011111" => data <= "110000";
        when "0111011100000000" => data <= "110000";
        when "0111011100000001" => data <= "110000";
        when "0111011100000010" => data <= "110000";
        when "0111011100000011" => data <= "110000";
        when "0111011100000100" => data <= "110000";
        when "0111011100000101" => data <= "110000";
        when "0111011100000110" => data <= "110000";
        when "0111011100000111" => data <= "110000";
        when "0111011100001000" => data <= "110000";
        when "0111011100001001" => data <= "110000";
        when "0111011100001010" => data <= "110000";
        when "0111011100001011" => data <= "110000";
        when "0111011100001100" => data <= "110000";
        when "0111011100001101" => data <= "110000";
        when "0111011100001110" => data <= "110000";
        when "0111011100001111" => data <= "110000";
        when "0111011100010000" => data <= "110000";
        when "0111011100010001" => data <= "110000";
        when "0111011100010010" => data <= "110000";
        when "0111011100010011" => data <= "110000";
        when "0111011100010100" => data <= "110000";
        when "0111011100010101" => data <= "110000";
        when "0111011100010110" => data <= "110000";
        when "0111011100010111" => data <= "110000";
        when "0111011100011000" => data <= "110000";
        when "0111011100011001" => data <= "110000";
        when "0111011100011010" => data <= "110000";
        when "0111011100011011" => data <= "110000";
        when "0111011100011100" => data <= "110000";
        when "0111011100011101" => data <= "110000";
        when "0111011100011110" => data <= "110000";
        when "0111011100011111" => data <= "110000";
        when "0111011100100000" => data <= "110000";
        when "0111011100100001" => data <= "110000";
        when "0111011100100010" => data <= "110000";
        when "0111011100100011" => data <= "110000";
        when "0111011100100100" => data <= "110000";
        when "0111011100100101" => data <= "110000";
        when "0111011100100110" => data <= "110000";
        when "0111011100100111" => data <= "110000";
        when "0111011100101000" => data <= "110000";
        when "0111011100101001" => data <= "110000";
        when "0111011100101010" => data <= "110000";
        when "0111011100101011" => data <= "110000";
        when "0111011100101100" => data <= "110000";
        when "0111011100101101" => data <= "110000";
        when "0111011100101110" => data <= "110000";
        when "0111011100101111" => data <= "110000";
        when "0111011100110000" => data <= "110000";
        when "0111011100110001" => data <= "110000";
        when "0111011100110010" => data <= "110000";
        when "0111011100110011" => data <= "110000";
        when "0111011100110100" => data <= "110000";
        when "0111011100110101" => data <= "110000";
        when "0111011100110110" => data <= "110000";
        when "0111011100110111" => data <= "110000";
        when "0111011100111000" => data <= "110000";
        when "0111011100111001" => data <= "110000";
        when "0111011100111010" => data <= "110000";
        when "0111011100111011" => data <= "110000";
        when "0111011100111100" => data <= "110000";
        when "0111011100111101" => data <= "110000";
        when "0111011100111110" => data <= "110000";
        when "0111011100111111" => data <= "110000";
        when "0111011101000000" => data <= "110000";
        when "0111011101000001" => data <= "110000";
        when "0111011101000010" => data <= "110000";
        when "0111011101000011" => data <= "110000";
        when "0111011101000100" => data <= "110000";
        when "0111011101000101" => data <= "110000";
        when "0111011101000110" => data <= "110000";
        when "0111011101000111" => data <= "110000";
        when "0111011101001000" => data <= "110000";
        when "0111011101001001" => data <= "110000";
        when "0111011101001010" => data <= "110000";
        when "0111011101001011" => data <= "110000";
        when "0111011101001100" => data <= "110000";
        when "0111011101001101" => data <= "110000";
        when "0111011101001110" => data <= "110000";
        when "0111011101001111" => data <= "110000";
        when "0111011101010000" => data <= "110000";
        when "0111011101010001" => data <= "110000";
        when "0111011101010010" => data <= "110000";
        when "0111011101010011" => data <= "110000";
        when "0111011101010100" => data <= "110000";
        when "0111011101010101" => data <= "110000";
        when "0111011101010110" => data <= "110000";
        when "0111011101010111" => data <= "110000";
        when "0111011101011000" => data <= "110000";
        when "0111011101011001" => data <= "110000";
        when "0111011101011010" => data <= "110000";
        when "0111011101011011" => data <= "110000";
        when "0111011101011100" => data <= "110000";
        when "0111011101011101" => data <= "110000";
        when "0111011101011110" => data <= "110000";
        when "0111011101011111" => data <= "110000";
        when "0111011101100000" => data <= "110000";
        when "0111011101100001" => data <= "110000";
        when "0111011101100010" => data <= "110000";
        when "0111011101100011" => data <= "110000";
        when "0111011101100100" => data <= "110000";
        when "0111011101100101" => data <= "110000";
        when "0111011101100110" => data <= "110000";
        when "0111011101100111" => data <= "110000";
        when "0111011101101000" => data <= "110000";
        when "0111011101101001" => data <= "110000";
        when "0111011101101010" => data <= "110000";
        when "0111011101101011" => data <= "110000";
        when "0111011101101100" => data <= "110000";
        when "0111011101101101" => data <= "110000";
        when "0111011101101110" => data <= "110000";
        when "0111011101101111" => data <= "110000";
        when "0111011101110000" => data <= "110000";
        when "0111011101110001" => data <= "110000";
        when "0111011101110010" => data <= "110000";
        when "0111011101110011" => data <= "110000";
        when "0111011101110100" => data <= "110000";
        when "0111011101110101" => data <= "110000";
        when "0111011101110110" => data <= "110000";
        when "0111011101110111" => data <= "110000";
        when "0111011101111000" => data <= "110000";
        when "0111011101111001" => data <= "110000";
        when "0111011101111010" => data <= "110000";
        when "0111011101111011" => data <= "110000";
        when "0111011101111100" => data <= "110000";
        when "0111011101111101" => data <= "110000";
        when "0111011101111110" => data <= "110000";
        when "0111011101111111" => data <= "110000";
        when "0111011110000000" => data <= "110000";
        when "0111011110000001" => data <= "110000";
        when "0111011110000010" => data <= "110000";
        when "0111011110000011" => data <= "110000";
        when "0111011110000100" => data <= "110000";
        when "0111011110000101" => data <= "110000";
        when "0111011110000110" => data <= "110000";
        when "0111011110000111" => data <= "110000";
        when "0111011110001000" => data <= "110000";
        when "0111011110001001" => data <= "110000";
        when "0111011110001010" => data <= "110000";
        when "0111011110001011" => data <= "110000";
        when "0111011110001100" => data <= "110000";
        when "0111011110001101" => data <= "110000";
        when "0111011110001110" => data <= "110000";
        when "0111011110001111" => data <= "110000";
        when "0111011110010000" => data <= "110000";
        when "0111011110010001" => data <= "110000";
        when "0111011110010010" => data <= "110000";
        when "0111011110010011" => data <= "110000";
        when "0111011110010100" => data <= "110000";
        when "0111011110010101" => data <= "110000";
        when "0111011110010110" => data <= "110000";
        when "0111011110010111" => data <= "110000";
        when "0111011110011000" => data <= "110000";
        when "0111011110011001" => data <= "110000";
        when "0111011110011010" => data <= "110000";
        when "0111011110011011" => data <= "110000";
        when "0111011110011100" => data <= "110000";
        when "0111011110011101" => data <= "110000";
        when "0111011110011110" => data <= "110000";
        when "0111011110011111" => data <= "110000";
        when others => data <= "000000";
      end case;
    end if;
  end process;
end;
